wbs_we_i
wbs_stb_i
wbs_sel_i_3_
wbs_sel_i_2_
wbs_sel_i_1_
wbs_sel_i_0_
wbs_rty_o
wbs_err_o
wbs_dat_o_9_
wbs_dat_o_8_
wbs_dat_o_7_
wbs_dat_o_6_
wbs_dat_o_5_
wbs_dat_o_4_
wbs_dat_o_3_
wbs_dat_o_31_
wbs_dat_o_30_
wbs_dat_o_2_
wbs_dat_o_29_
wbs_dat_o_28_
wbs_dat_o_27_
wbs_dat_o_26_
wbs_dat_o_25_
wbs_dat_o_24_
wbs_dat_o_23_
wbs_dat_o_22_
wbs_dat_o_21_
wbs_dat_o_20_
wbs_dat_o_1_
wbs_dat_o_19_
wbs_dat_o_18_
wbs_dat_o_17_
wbs_dat_o_16_
wbs_dat_o_15_
wbs_dat_o_14_
wbs_dat_o_13_
wbs_dat_o_12_
wbs_dat_o_11_
wbs_dat_o_10_
wbs_dat_o_0_
wbs_dat_i_9_
wbs_dat_i_8_
wbs_dat_i_7_
wbs_dat_i_6_
wbs_dat_i_5_
wbs_dat_i_4_
wbs_dat_i_3_
wbs_dat_i_31_
wbs_dat_i_30_
wbs_dat_i_2_
wbs_dat_i_29_
wbs_dat_i_28_
wbs_dat_i_27_
wbs_dat_i_26_
wbs_dat_i_25_
wbs_dat_i_24_
wbs_dat_i_23_
wbs_dat_i_22_
wbs_dat_i_21_
wbs_dat_i_20_
wbs_dat_i_1_
wbs_dat_i_19_
wbs_dat_i_18_
wbs_dat_i_17_
wbs_dat_i_16_
wbs_dat_i_15_
wbs_dat_i_14_
wbs_dat_i_13_
wbs_dat_i_12_
wbs_dat_i_11_
wbs_dat_i_10_
wbs_dat_i_0_
wbs_cyc_i
wbs_cti_i_2_
wbs_cti_i_1_
wbs_cti_i_0_
wbs_bte_i_1_
wbs_bte_i_0_
wbs_adr_i_9_
wbs_adr_i_8_
wbs_adr_i_7_
wbs_adr_i_6_
wbs_adr_i_5_
wbs_adr_i_4_
wbs_adr_i_3_
wbs_adr_i_31_
wbs_adr_i_30_
wbs_adr_i_2_
wbs_adr_i_29_
wbs_adr_i_28_
wbs_adr_i_27_
wbs_adr_i_26_
wbs_adr_i_25_
wbs_adr_i_24_
wbs_adr_i_23_
wbs_adr_i_22_
wbs_adr_i_21_
wbs_adr_i_20_
wbs_adr_i_1_
wbs_adr_i_19_
wbs_adr_i_18_
wbs_adr_i_17_
wbs_adr_i_16_
wbs_adr_i_15_
wbs_adr_i_14_
wbs_adr_i_13_
wbs_adr_i_12_
wbs_adr_i_11_
wbs_adr_i_10_
wbs_adr_i_0_
wbs_ack_o
wbm_we_o
wbm_stb_o
wbm_sel_o_3_
wbm_sel_o_2_
wbm_sel_o_1_
wbm_sel_o_0_
wbm_rty_i
wbm_err_i
wbm_dat_o_9_
wbm_dat_o_8_
wbm_dat_o_7_
wbm_dat_o_6_
wbm_dat_o_5_
wbm_dat_o_4_
wbm_dat_o_3_
wbm_dat_o_31_
wbm_dat_o_30_
wbm_dat_o_2_
wbm_dat_o_29_
wbm_dat_o_28_
wbm_dat_o_27_
wbm_dat_o_26_
wbm_dat_o_25_
wbm_dat_o_24_
wbm_dat_o_23_
wbm_dat_o_22_
wbm_dat_o_21_
wbm_dat_o_20_
wbm_dat_o_1_
wbm_dat_o_19_
wbm_dat_o_18_
wbm_dat_o_17_
wbm_dat_o_16_
wbm_dat_o_15_
wbm_dat_o_14_
wbm_dat_o_13_
wbm_dat_o_12_
wbm_dat_o_11_
wbm_dat_o_10_
wbm_dat_o_0_
wbm_dat_i_9_
wbm_dat_i_8_
wbm_dat_i_7_
wbm_dat_i_6_
wbm_dat_i_5_
wbm_dat_i_4_
wbm_dat_i_3_
wbm_dat_i_31_
wbm_dat_i_30_
wbm_dat_i_2_
wbm_dat_i_29_
wbm_dat_i_28_
wbm_dat_i_27_
wbm_dat_i_26_
wbm_dat_i_25_
wbm_dat_i_24_
wbm_dat_i_23_
wbm_dat_i_22_
wbm_dat_i_21_
wbm_dat_i_20_
wbm_dat_i_1_
wbm_dat_i_19_
wbm_dat_i_18_
wbm_dat_i_17_
wbm_dat_i_16_
wbm_dat_i_15_
wbm_dat_i_14_
wbm_dat_i_13_
wbm_dat_i_12_
wbm_dat_i_11_
wbm_dat_i_10_
wbm_dat_i_0_
wbm_cyc_o
wbm_cti_o_2_
wbm_cti_o_1_
wbm_cti_o_0_
wbm_adr_o_9_
wbm_adr_o_8_
wbm_adr_o_7_
wbm_adr_o_6_
wbm_adr_o_5_
wbm_adr_o_4_
wbm_adr_o_3_
wbm_adr_o_31_
wbm_adr_o_30_
wbm_adr_o_2_
wbm_adr_o_29_
wbm_adr_o_28_
wbm_adr_o_27_
wbm_adr_o_26_
wbm_adr_o_25_
wbm_adr_o_24_
wbm_adr_o_23_
wbm_adr_o_22_
wbm_adr_o_21_
wbm_adr_o_20_
wbm_adr_o_1_
wbm_adr_o_19_
wbm_adr_o_18_
wbm_adr_o_17_
wbm_adr_o_16_
wbm_adr_o_15_
wbm_adr_o_14_
wbm_adr_o_13_
wbm_adr_o_12_
wbm_adr_o_11_
wbm_adr_o_10_
wbm_adr_o_0_
wbm_ack_i
wb_rst_o
wb_int_i
pci_trdy_oe_o
pci_trdy_o
pci_trdy_i
pci_stop_oe_o
pci_stop_o
pci_stop_i
pci_serr_oe_o
pci_serr_o
pci_rst_oe_o
pci_rst_i
pci_req_oe_o
pci_req_o
pci_perr_oe_o
pci_perr_o
pci_perr_i
pci_par_oe_o
pci_par_o
pci_par_i
pci_irdy_oe_o
pci_irdy_o
pci_irdy_i
pci_inta_oe_o
pci_idsel_i
pci_gnt_i
pci_frame_oe_o
pci_frame_o
pci_frame_i
pci_devsel_oe_o
pci_devsel_o
pci_devsel_i
pci_cbe_oe_o_3_
pci_cbe_oe_o_2_
pci_cbe_oe_o_1_
pci_cbe_oe_o_0_
pci_cbe_o_3_
pci_cbe_o_2_
pci_cbe_o_1_
pci_cbe_o_0_
pci_cbe_i_3_
pci_cbe_i_2_
pci_cbe_i_1_
pci_cbe_i_0_
pci_ad_oe_o_9_
pci_ad_oe_o_8_
pci_ad_oe_o_7_
pci_ad_oe_o_6_
pci_ad_oe_o_5_
pci_ad_oe_o_4_
pci_ad_oe_o_3_
pci_ad_oe_o_31_
pci_ad_oe_o_30_
pci_ad_oe_o_2_
pci_ad_oe_o_29_
pci_ad_oe_o_28_
pci_ad_oe_o_27_
pci_ad_oe_o_26_
pci_ad_oe_o_25_
pci_ad_oe_o_24_
pci_ad_oe_o_23_
pci_ad_oe_o_22_
pci_ad_oe_o_21_
pci_ad_oe_o_20_
pci_ad_oe_o_1_
pci_ad_oe_o_19_
pci_ad_oe_o_18_
pci_ad_oe_o_17_
pci_ad_oe_o_16_
pci_ad_oe_o_15_
pci_ad_oe_o_14_
pci_ad_oe_o_13_
pci_ad_oe_o_12_
pci_ad_oe_o_11_
pci_ad_oe_o_10_
pci_ad_oe_o_0_
pci_ad_o_9_
pci_ad_o_8_
pci_ad_o_7_
pci_ad_o_6_
pci_ad_o_5_
pci_ad_o_4_
pci_ad_o_3_
pci_ad_o_31_
pci_ad_o_30_
pci_ad_o_2_
pci_ad_o_29_
pci_ad_o_28_
pci_ad_o_27_
pci_ad_o_26_
pci_ad_o_25_
pci_ad_o_24_
pci_ad_o_23_
pci_ad_o_22_
pci_ad_o_21_
pci_ad_o_20_
pci_ad_o_1_
pci_ad_o_19_
pci_ad_o_18_
pci_ad_o_17_
pci_ad_o_16_
pci_ad_o_15_
pci_ad_o_14_
pci_ad_o_13_
pci_ad_o_12_
pci_ad_o_11_
pci_ad_o_10_
pci_ad_o_0_
pci_ad_i_9_
pci_ad_i_8_
pci_ad_i_7_
pci_ad_i_6_
pci_ad_i_5_
pci_ad_i_4_
pci_ad_i_3_
pci_ad_i_31_
pci_ad_i_30_
pci_ad_i_2_
pci_ad_i_29_
pci_ad_i_28_
pci_ad_i_27_
pci_ad_i_26_
pci_ad_i_25_
pci_ad_i_24_
pci_ad_i_23_
pci_ad_i_22_
pci_ad_i_21_
pci_ad_i_20_
pci_ad_i_1_
pci_ad_i_19_
pci_ad_i_18_
pci_ad_i_17_
pci_ad_i_16_
pci_ad_i_15_
pci_ad_i_14_
pci_ad_i_13_
pci_ad_i_12_
pci_ad_i_11_
pci_ad_i_10_
pci_ad_i_0_
FE_OCPN1849_n_16798
FE_OCPN1850_n_16486
FE_OCPN1851_n_16486
FE_OCPN1852_n_14981
FE_OCPN1853_n_14981
FE_OCPN1854_n_16949
FE_OCPN1855_n_16949
FE_OCPN1856_n_12030
FE_OCPN1857_n_12030
FE_OCPN1860_n_14971
FE_OCPN1861_n_14971
FE_OCPN1862_n_15808
FE_OCPN1863_n_15808
FE_OCPN1864_n_15808
FE_OCPN1865_n_15808
FE_OCPN1866_n_15808
FE_OCPN1867_n_15768
FE_OCPN1868_n_15768
FE_OCPN1869_n_15371
FE_OCPN1870_n_15371
FE_OCPN1871_n_12099
FE_OCPN1872_n_12099
FE_OCPN1873_n_12099
FE_OCPN1874_FE_OFN1678_n_10588
FE_OCPN1875_FE_OFN1678_n_10588
FE_OCPN1876_n_15978
FE_OCPN1877_n_15978
FE_OCPN1879_n_9991
FE_OCPN1880_FE_OFN941_n_16089
FE_OCPN1881_FE_OFN941_n_16089
FE_OCPN1884_FE_OFN1454_n_12028
FE_OCPN1885_FE_OFN1454_n_12028
FE_OCPN1888_n_12357
FE_OCPN1889_n_12357
FE_OCPN1890_FE_OFN1430_n_12104
FE_OCPN1891_FE_OFN1430_n_12104
FE_OCPN1894_parchk_pci_ad_reg_in_1228
FE_OCPN1895_parchk_pci_ad_reg_in_1228
FE_OCPN1896_parchk_pci_ad_reg_in_1228
FE_OCPN1897_parchk_pci_ad_reg_in_1228
FE_OCPN1898_n_1061
FE_OCPN1899_n_1061
FE_OCPN1900_n_2071
FE_OCPN1901_n_2071
FE_OCPN1902_FE_OFN1677_n_10588
FE_OCPN1903_FE_OFN1677_n_10588
FE_OCPN1904_n_11884
FE_OCPN1905_n_11884
FE_OCPN1906_FE_OFN1754_n_12681
FE_OCPN1907_FE_OFN1754_n_12681
FE_OCPN1908_parchk_pci_ad_reg_in_1231
FE_OCPN1909_parchk_pci_ad_reg_in_1231
FE_OCPN1910_parchk_pci_ad_reg_in_1231
FE_OCPN1911_parchk_pci_ad_reg_in_1229
FE_OCPN1912_parchk_pci_ad_reg_in_1229
FE_OCPN1913_parchk_pci_ad_reg_in_1229
FE_OCPN1914_parchk_pci_ad_reg_in_1229
FE_OCPN1915_n_16289
FE_OCPN1916_n_16289
FE_OCPN1917_n_1291
FE_OCPN1918_n_1291
FE_OCPN1919_n_8927
FE_OCPN1920_n_8927
FE_OCPN1921_n_8927
FE_OCPN1922_FE_OFN1685_n_16891
FE_OCPN1923_FE_OFN1685_n_16891
FE_OCPN1925_FE_OFN1758_n_13997
FE_OCPN1927_n_7102
FE_OCPN1928_parchk_pci_ad_reg_in_1226
FE_OCPN1929_parchk_pci_ad_reg_in_1226
FE_OCPN1930_parchk_pci_ad_reg_in_1226
FE_OCPN1931_parchk_pci_ad_reg_in_1226
FE_OCPN1932_FE_OFN1697_n_9975
FE_OCPN1933_FE_OFN1697_n_9975
FE_OCPN1936_n_15566
FE_OCPN1937_FE_OFN1683_n_16891
FE_OCPN1938_FE_OFN1683_n_16891
FE_OCPN1941_n_11823
FE_OCPN1942_n_11823
FE_OCPN1943_FE_OFN1731_n_11019
FE_OCPN1944_FE_OFN1731_n_11019
FE_OCPN1945_FE_OFN130_n_12104
FE_OCPN1946_FE_OFN130_n_12104
FE_OCPN1947_FE_OFN1430_n_12104
FE_OCPN1948_FE_OFN1430_n_12104
FE_OCPN1950_n_12030
FE_OCPN1951_FE_OFN1753_n_12681
FE_OCPN1952_FE_OFN1753_n_12681
FE_OCPN1953_parchk_pci_ad_reg_in_1225
FE_OCPN1954_parchk_pci_ad_reg_in_1225
FE_OCPN1955_parchk_pci_ad_reg_in_1225
FE_OCPN1956_parchk_pci_ad_reg_in_1225
FE_OCPN1957_FE_OFN119_n_12502
FE_OCPN1958_FE_OFN119_n_12502
FE_OCPN1959_n_16495
FE_OCPN1960_n_16495
FE_OCPN1961_n_16495
FE_OCPN1962_parchk_pci_ad_reg_in_1227
FE_OCPN1963_parchk_pci_ad_reg_in_1227
FE_OCPN1964_parchk_pci_ad_reg_in_1227
FE_OCPN1965_parchk_pci_ad_reg_in_1227
FE_OCPN1970_n_15445
FE_OCPN1971_n_15445
FE_OCPN1972_n_3252
FE_OCPN1973_n_3252
FE_OCPN1975_FE_OFN961_n_16810
FE_OCPN1976_FE_OFN1367_n_15587
FE_OCPN1977_FE_OFN1367_n_15587
FE_OCPN1978_FE_OFN1722_n_16317
FE_OCPN1979_FE_OFN1722_n_16317
FE_OCPN1980_FE_OFN1719_n_16317
FE_OCPN1981_FE_OFN1719_n_16317
FE_OCPN1986_n_7102
FE_OCPN1987_FE_OFN1264_n_8567
FE_OCPN1988_FE_OFN1264_n_8567
FE_OCPN1990_n_16000
FE_OCPN1991_n_16000
FE_OCPN1992_g66358_p
FE_OCPN1993_g66358_p
FE_OCPN1995_n_9991
FE_OCPN1997_FE_OFN1711_n_9320
FE_OCPN1998_n_13743
FE_OCPN1999_n_13743
FE_OCPN2000_n_13743
FE_OCPN2001_n_11884
FE_OCPN2002_n_11884
FE_OCPN2004_n_11823
FE_OCPN2020_parchk_pci_ad_reg_in_1222
FE_OCPN2021_parchk_pci_ad_reg_in_1222
FE_OCPN2022_parchk_pci_ad_reg_in_1222
FE_OCPN2029_n_10763
FE_OCPN2030_n_10763
FE_OCPN2042_FE_OFN675_n_8140
FE_OCPN2043_FE_OFN675_n_8140
FE_OCPN2119_FE_OFN448_n_10853
FE_OCPN2120_FE_OFN448_n_10853
FE_OCPUNCON2033_n_14837
FE_OCPUNCON2034_n_14837
FE_OCP_DRV_N2035_n_1805
FE_OCP_DRV_N2036_n_1805
FE_OCP_DRV_N2040_n_8660
FE_OCP_DRV_N2041_n_8660
FE_OCP_RBN1982_n_15919
FE_OCP_RBN1983_n_15919
FE_OCP_RBN1984_n_15919
FE_OCP_RBN2005_wbs_cti_i_1_
FE_OCP_RBN2006_n_16523
FE_OCP_RBN2007_n_16523
FE_OCP_RBN2008_FE_RN_290_0
FE_OCP_RBN2010_FE_RN_290_0
FE_OCP_RBN2011_FE_OFN1725_n_14987
FE_OCP_RBN2031_n_10244
FE_OCP_RBN2032_n_10244
FE_OCP_RBN2037_FE_OCPN2000_n_13743
FE_OCP_RBN2038_FE_OCPN2000_n_13743
FE_OCP_RBN2039_FE_OCPN2000_n_13743
FE_OCP_RBN2044_n_16533
FE_OCP_RBN2045_n_16533
FE_OCP_RBN2046_n_16533
FE_OCP_RBN2055_FE_RN_356_0
FE_OCP_RBN2056_FE_RN_356_0
FE_OCP_RBN2057_FE_RN_378_0
FE_OCP_RBN2058_FE_RN_378_0
FE_OCP_RBN2059_FE_RN_378_0
FE_OCP_RBN2060_FE_RN_378_0
FE_OCP_RBN2061_FE_RN_378_0
FE_OCP_RBN2062_n_16572
FE_OCP_RBN2063_n_16572
FE_OCP_RBN2064_n_16572
FE_OCP_RBN2065_n_16572
FE_OCP_RBN2069_n_16572
FE_OCP_RBN2071_n_9155
FE_OCP_RBN2074_n_11767
FE_OCP_RBN2076_n_11767
FE_OCP_RBN2077_n_16975
FE_OCP_RBN2080_n_16975
FE_OCP_RBN2081_n_16975
FE_OCP_RBN2082_n_10244
FE_OCP_RBN2084_n_10244
FE_OCP_RBN2085_FE_OFN1756_n_13997
FE_OCP_RBN2086_FE_OFN1756_n_13997
FE_OCP_RBN2087_FE_OFN1756_n_13997
FE_OCP_RBN2089_FE_OFN1433_n_12042
FE_OCP_RBN2091_FE_OFN1746_n_11027
FE_OCP_RBN2092_FE_OFN1746_n_11027
FE_OCP_RBN2093_FE_OFN1746_n_11027
FE_OCP_RBN2094_FE_OCPN1856_n_12030
FE_OCP_RBN2095_FE_OCPN1856_n_12030
FE_OCP_RBN2099_pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_1_
FE_OCP_RBN2100_n_15347
FE_OCP_RBN2101_n_15347
FE_OCP_RBN2102_FE_RN_255_0
FE_OCP_RBN2103_FE_RN_255_0
FE_OCP_RBN2104_n_9155
FE_OCP_RBN2105_n_9155
FE_OCP_RBN2106_n_9155
FE_OCP_RBN2107_n_9155
FE_OCP_RBN2108_n_8872
FE_OCP_RBN2109_n_8872
FE_OCP_RBN2110_n_8872
FE_OCP_RBN2111_n_8872
FE_OCP_RBN2112_n_8872
FE_OCP_RBN2113_n_8872
FE_OCP_RBN2115_n_16553
FE_OCP_RBN2116_n_16553
FE_OCP_RBN2117_n_16553
FE_OCP_RBN2118_n_16553
FE_OCP_RBN2121_n_16966
FE_OCP_RBN2122_n_16966
FE_OCP_RBN2123_n_16966
FE_OCP_RBN2124_n_16966
FE_OFN1000_n_7350
FE_OFN1004_n_13221
FE_OFN1005_n_13221
FE_OFN1006_n_13221
FE_OFN1007_n_13221
FE_OFN1008_n_13221
FE_OFN1009_n_13221
FE_OFN1010_g64577_p
FE_OFN1011_g64577_p
FE_OFN1012_g64577_p
FE_OFN1013_g64577_p
FE_OFN1015_g64577_p
FE_OFN1016_g64577_p
FE_OFN1017_g64577_p
FE_OFN1018_g64577_p
FE_OFN1019_g64577_p
FE_OFN1022_g64577_p
FE_OFN1023_g64577_p
FE_OFN1024_g64577_p
FE_OFN1026_g64577_p
FE_OFN1027_g64577_p
FE_OFN1028_g64577_p
FE_OFN1029_g64577_p
FE_OFN1032_g64577_p
FE_OFN1033_g64577_p
FE_OFN1034_g64577_p
FE_OFN1035_g64577_p
FE_OFN1038_g64577_p
FE_OFN1040_g64577_p
FE_OFN1041_g64577_p
FE_OFN1042_g64577_p
FE_OFN1043_g64577_p
FE_OFN1046_g64577_p
FE_OFN1047_g64577_p
FE_OFN1048_g64577_p
FE_OFN1050_g64577_p
FE_OFN1051_g64577_p
FE_OFN1052_g64577_p
FE_OFN1054_g64577_p
FE_OFN1055_g64577_p
FE_OFN1057_g64577_p
FE_OFN1058_g64577_p
FE_OFN1059_g64577_p
FE_OFN1062_n_8176
FE_OFN1063_n_8176
FE_OFN1064_n_8176
FE_OFN1065_n_8176
FE_OFN1066_n_8176
FE_OFN1067_n_8176
FE_OFN1068_n_8176
FE_OFN1069_n_8069
FE_OFN1070_n_8069
FE_OFN1071_n_8069
FE_OFN1072_n_8069
FE_OFN1073_n_8069
FE_OFN1074_n_7845
FE_OFN1075_n_7845
FE_OFN1076_n_7845
FE_OFN1077_n_7845
FE_OFN1078_n_7845
FE_OFN1079_n_7845
FE_OFN1080_n_13249
FE_OFN1081_n_13249
FE_OFN1082_n_13249
FE_OFN1083_n_13249
FE_OFN1084_n_13249
FE_OFN1085_n_13249
FE_OFN1087_n_15325
FE_OFN1088_n_15325
FE_OFN1089_n_15325
FE_OFN108_n_12028
FE_OFN1090_n_5615
FE_OFN1091_n_5615
FE_OFN1092_n_5615
FE_OFN1093_n_5615
FE_OFN1094_n_5615
FE_OFN1095_n_5592
FE_OFN1099_n_5592
FE_OFN10_n_11877
FE_OFN1100_n_5592
FE_OFN1101_n_5592
FE_OFN1103_n_5592
FE_OFN1105_n_3476
FE_OFN1106_n_3476
FE_OFN1107_n_3476
FE_OFN1108_n_3476
FE_OFN1109_n_3476
FE_OFN1110_n_3476
FE_OFN1111_n_3476
FE_OFN1112_n_3476
FE_OFN1113_n_3476
FE_OFN1114_n_3476
FE_OFN1115_n_5742
FE_OFN1116_n_5742
FE_OFN1117_n_5742
FE_OFN1118_n_6935
FE_OFN1119_n_6935
FE_OFN1120_n_6935
FE_OFN1123_n_6935
FE_OFN1124_n_6935
FE_OFN1125_n_4090
FE_OFN1126_n_4090
FE_OFN1127_n_4090
FE_OFN1128_n_4090
FE_OFN1129_n_4090
FE_OFN1130_n_6356
FE_OFN1131_n_6356
FE_OFN1132_n_6356
FE_OFN1133_n_6356
FE_OFN1134_n_4151
FE_OFN1135_n_4151
FE_OFN1136_n_4151
FE_OFN1137_n_4151
FE_OFN1138_n_4151
FE_OFN1139_n_6886
FE_OFN1140_n_6886
FE_OFN1141_n_6886
FE_OFN1143_n_6391
FE_OFN1146_n_6391
FE_OFN1147_n_6391
FE_OFN1148_n_6391
FE_OFN1149_n_6391
FE_OFN1150_n_6391
FE_OFN1151_n_6391
FE_OFN1152_n_6391
FE_OFN1156_n_6391
FE_OFN1157_n_6391
FE_OFN1159_n_6391
FE_OFN1160_n_6391
FE_OFN1161_n_6391
FE_OFN1162_n_6391
FE_OFN1163_n_4092
FE_OFN1164_n_4092
FE_OFN1165_n_4092
FE_OFN1166_n_4092
FE_OFN1167_n_4092
FE_OFN1168_n_4093
FE_OFN1169_n_4093
FE_OFN1170_n_4093
FE_OFN1173_n_4093
FE_OFN1174_n_4093
FE_OFN1175_n_4093
FE_OFN1176_n_4093
FE_OFN1177_n_4143
FE_OFN117_n_12306
FE_OFN1181_n_4143
FE_OFN1182_n_4143
FE_OFN1184_n_4143
FE_OFN1185_n_4143
FE_OFN1186_n_4095
FE_OFN1187_n_4095
FE_OFN1188_n_4095
FE_OFN1189_n_4095
FE_OFN1190_n_4095
FE_OFN1191_n_4095
FE_OFN1192_n_4095
FE_OFN1193_n_4095
FE_OFN1194_n_4096
FE_OFN1195_n_4096
FE_OFN1196_n_4096
FE_OFN1197_n_4096
FE_OFN1198_n_4096
FE_OFN1199_n_4096
FE_OFN119_n_12502
FE_OFN11_n_11877
FE_OFN1204_n_4097
FE_OFN1205_n_4097
FE_OFN1206_n_4097
FE_OFN1207_n_4097
FE_OFN1208_n_4098
FE_OFN1209_n_4098
FE_OFN1210_n_4098
FE_OFN1211_n_4098
FE_OFN1212_n_4098
FE_OFN1213_n_4098
FE_OFN1214_n_5763
FE_OFN1215_n_5763
FE_OFN1216_n_5763
FE_OFN1217_n_5763
FE_OFN1218_n_5763
FE_OFN1219_n_13124
FE_OFN1220_n_13124
FE_OFN1221_n_13124
FE_OFN1222_n_13124
FE_OFN1223_n_6624
FE_OFN1225_n_6624
FE_OFN1226_n_6624
FE_OFN1227_n_6624
FE_OFN1229_n_6624
FE_OFN1231_n_6624
FE_OFN1232_n_6624
FE_OFN1233_n_6624
FE_OFN1234_n_6624
FE_OFN1235_n_6436
FE_OFN1236_n_6436
FE_OFN1237_n_6436
FE_OFN1238_n_6436
FE_OFN1239_n_6436
FE_OFN1241_n_13668
FE_OFN1242_n_13652
FE_OFN1243_n_13652
FE_OFN1244_n_13560
FE_OFN1245_n_13560
FE_OFN1246_n_13671
FE_OFN1247_n_13671
FE_OFN1248_n_16439
FE_OFN1249_n_16439
FE_OFN1250_n_16439
FE_OFN1251_n_16439
FE_OFN1252_n_16439
FE_OFN1253_n_8567
FE_OFN1254_n_8567
FE_OFN1255_n_8567
FE_OFN1257_n_8567
FE_OFN1258_n_8567
FE_OFN1259_n_8567
FE_OFN1260_n_8567
FE_OFN1261_n_8567
FE_OFN1262_n_8567
FE_OFN1263_n_8567
FE_OFN1264_n_8567
FE_OFN1265_n_8567
FE_OFN1266_n_8567
FE_OFN1267_n_8567
FE_OFN1268_n_8567
FE_OFN1269_n_8567
FE_OFN1270_n_8567
FE_OFN1271_n_8567
FE_OFN1272_n_8567
FE_OFN1273_n_8567
FE_OFN1274_n_8567
FE_OFN1275_n_8567
FE_OFN1276_n_8567
FE_OFN1277_n_8567
FE_OFN1279_n_8567
FE_OFN1280_n_8567
FE_OFN1281_n_8567
FE_OFN1282_n_8567
FE_OFN1283_n_8567
FE_OFN1284_n_8567
FE_OFN1285_n_8567
FE_OFN1286_n_8567
FE_OFN1287_n_8567
FE_OFN1288_n_8567
FE_OFN1289_n_8567
FE_OFN1290_n_8567
FE_OFN1291_n_8567
FE_OFN1292_n_8567
FE_OFN1293_n_8567
FE_OFN1294_n_8567
FE_OFN1295_n_8567
FE_OFN1296_n_8567
FE_OFN1297_n_8567
FE_OFN1298_n_8567
FE_OFN1299_n_8567
FE_OFN129_n_12104
FE_OFN12_n_11877
FE_OFN1300_n_8567
FE_OFN1301_n_8567
FE_OFN1302_n_8567
FE_OFN1303_n_8567
FE_OFN1304_n_8567
FE_OFN1305_n_8567
FE_OFN1306_n_8567
FE_OFN1307_n_8567
FE_OFN1308_n_8567
FE_OFN1309_n_8567
FE_OFN130_n_12104
FE_OFN1310_n_8567
FE_OFN1311_n_8567
FE_OFN1312_n_8567
FE_OFN1313_n_8567
FE_OFN1314_n_8567
FE_OFN1315_n_8567
FE_OFN1316_n_8567
FE_OFN1317_n_8567
FE_OFN1318_n_8567
FE_OFN1319_n_8567
FE_OFN1320_n_8567
FE_OFN1321_n_8567
FE_OFN1322_n_8567
FE_OFN1323_n_8567
FE_OFN1324_n_16779
FE_OFN1325_n_16779
FE_OFN1326_n_16779
FE_OFN1327_n_16779
FE_OFN1328_n_16301
FE_OFN1329_n_16301
FE_OFN1330_n_16301
FE_OFN1331_n_16301
FE_OFN1332_n_16301
FE_OFN1334_n_9372
FE_OFN1336_n_9372
FE_OFN1337_n_9372
FE_OFN1338_n_9372
FE_OFN1339_n_9372
FE_OFN1340_n_9372
FE_OFN1341_n_9372
FE_OFN1342_n_11125
FE_OFN1343_n_11125
FE_OFN1344_n_11125
FE_OFN1345_n_11125
FE_OFN1346_n_11125
FE_OFN1347_n_11125
FE_OFN1348_n_9163
FE_OFN1349_n_9163
FE_OFN1350_n_15558
FE_OFN1351_n_15558
FE_OFN1352_n_15558
FE_OFN1353_n_15558
FE_OFN1354_n_15558
FE_OFN1355_n_15558
FE_OFN1356_n_15558
FE_OFN1357_n_16698
FE_OFN1358_n_16698
FE_OFN1359_n_16698
FE_OFN1360_n_16698
FE_OFN1361_n_16698
FE_OFN1362_n_15587
FE_OFN1363_n_15587
FE_OFN1364_n_15587
FE_OFN1365_n_15587
FE_OFN1366_n_15587
FE_OFN1367_n_15587
FE_OFN1368_n_15587
FE_OFN1369_n_10538
FE_OFN1370_n_10538
FE_OFN1371_n_10538
FE_OFN1372_n_10538
FE_OFN1373_n_10538
FE_OFN1374_n_10853
FE_OFN1375_n_10853
FE_OFN1376_n_10853
FE_OFN1377_n_10853
FE_OFN1378_n_10853
FE_OFN1382_n_10143
FE_OFN1383_n_10143
FE_OFN1384_n_10143
FE_OFN1385_n_10143
FE_OFN1386_n_10143
FE_OFN1387_n_10143
FE_OFN1388_n_10143
FE_OFN1389_n_10595
FE_OFN1390_n_10595
FE_OFN1391_n_10595
FE_OFN1392_n_10595
FE_OFN1393_n_10595
FE_OFN1394_n_10566
FE_OFN1395_n_10566
FE_OFN1396_n_10566
FE_OFN1397_n_10566
FE_OFN1398_n_10566
FE_OFN1399_n_10566
FE_OFN13_n_11877
FE_OFN1400_n_10566
FE_OFN1401_n_11138
FE_OFN1402_n_11138
FE_OFN1403_n_11138
FE_OFN1404_n_11138
FE_OFN1405_n_11138
FE_OFN1406_n_11138
FE_OFN1407_n_11795
FE_OFN1408_n_11795
FE_OFN1409_n_11795
FE_OFN1411_n_11795
FE_OFN1412_n_11795
FE_OFN1413_n_11795
FE_OFN1414_n_10789
FE_OFN1415_n_10789
FE_OFN1416_n_10789
FE_OFN1417_n_10789
FE_OFN1418_n_10789
FE_OFN1419_g52675_p
FE_OFN1420_g52675_p
FE_OFN1421_g52675_p
FE_OFN1422_g52675_p
FE_OFN1423_g52675_p
FE_OFN1424_n_15768
FE_OFN1425_n_15768
FE_OFN1426_n_15768
FE_OFN1427_n_12104
FE_OFN1429_n_12104
FE_OFN1430_n_12104
FE_OFN1431_n_12104
FE_OFN1432_n_12042
FE_OFN1435_n_12042
FE_OFN1437_n_12042
FE_OFN1438_n_12042
FE_OFN1441_n_12502
FE_OFN1442_n_12502
FE_OFN1443_n_12502
FE_OFN1444_n_12502
FE_OFN1445_n_12502
FE_OFN1446_n_10780
FE_OFN1447_n_10780
FE_OFN1448_n_10780
FE_OFN1449_n_10780
FE_OFN1450_n_10780
FE_OFN1451_n_10780
FE_OFN1455_n_12028
FE_OFN1457_n_12306
FE_OFN1458_n_12306
FE_OFN1460_n_12306
FE_OFN1461_n_12306
FE_OFN1462_n_13736
FE_OFN1463_n_13736
FE_OFN1464_n_13736
FE_OFN1465_n_13736
FE_OFN1466_n_13736
FE_OFN1467_n_13741
FE_OFN1468_n_13741
FE_OFN1469_n_13741
FE_OFN1470_n_13741
FE_OFN1471_n_13741
FE_OFN1472_n_13741
FE_OFN1474_n_14995
FE_OFN1475_n_14995
FE_OFN1476_n_13995
FE_OFN1477_n_13995
FE_OFN1478_n_13995
FE_OFN1479_n_13995
FE_OFN1480_n_13995
FE_OFN1481_n_13995
FE_OFN1484_n_15366
FE_OFN1485_n_15366
FE_OFN1486_n_659
FE_OFN1488_n_15978
FE_OFN1489_n_15978
FE_OFN1490_n_15978
FE_OFN1491_n_1787
FE_OFN1492_n_1787
FE_OFN1493_n_1787
FE_OFN1494_n_1787
FE_OFN1495_n_1787
FE_OFN1496_n_9864
FE_OFN1497_n_9864
FE_OFN1498_n_9864
FE_OFN1499_n_9864
FE_OFN1500_n_9864
FE_OFN1501_n_9531
FE_OFN1502_n_9531
FE_OFN1503_n_9531
FE_OFN1504_n_9531
FE_OFN1505_n_9531
FE_OFN1506_n_9531
FE_OFN1507_n_4460
FE_OFN1508_n_4460
FE_OFN1509_n_4460
FE_OFN1510_n_4460
FE_OFN1511_n_4460
FE_OFN1512_n_4677
FE_OFN1513_n_4677
FE_OFN1514_n_4677
FE_OFN1515_n_4677
FE_OFN1516_n_4677
FE_OFN1517_n_4677
FE_OFN1518_n_4730
FE_OFN1519_n_4730
FE_OFN1520_n_4730
FE_OFN1521_n_4730
FE_OFN1522_n_4730
FE_OFN1523_n_4730
FE_OFN1524_n_4730
FE_OFN1525_n_4730
FE_OFN1527_n_4671
FE_OFN1529_n_4671
FE_OFN1530_n_4671
FE_OFN1531_n_4671
FE_OFN1532_n_4671
FE_OFN1533_n_9428
FE_OFN1534_n_9428
FE_OFN1535_n_9428
FE_OFN1536_n_9428
FE_OFN1537_n_9428
FE_OFN1538_n_9428
FE_OFN1539_n_9502
FE_OFN1540_n_9502
FE_OFN1541_n_9502
FE_OFN1542_n_9502
FE_OFN1543_n_9502
FE_OFN1544_n_9502
FE_OFN1545_n_4501
FE_OFN1546_n_4501
FE_OFN1547_n_4501
FE_OFN1548_n_4501
FE_OFN1549_n_4501
FE_OFN1550_n_4501
FE_OFN1552_n_4732
FE_OFN1553_n_4732
FE_OFN1554_n_4732
FE_OFN1555_n_4732
FE_OFN1556_n_4732
FE_OFN1557_n_4732
FE_OFN1558_n_4732
FE_OFN1559_n_4732
FE_OFN1560_n_2037
FE_OFN1561_n_2037
FE_OFN1562_n_2037
FE_OFN1563_n_2037
FE_OFN1564_n_9477
FE_OFN1565_n_9477
FE_OFN1566_n_9477
FE_OFN1567_n_9477
FE_OFN1568_n_9477
FE_OFN1569_n_9477
FE_OFN1570_n_9477
FE_OFN1571_n_9477
FE_OFN1572_n_9477
FE_OFN1573_n_9477
FE_OFN1574_n_9477
FE_OFN1575_n_9477
FE_OFN1578_n_16657
FE_OFN1579_n_16657
FE_OFN1580_n_16657
FE_OFN1581_n_16657
FE_OFN1582_n_16657
FE_OFN1583_n_16657
FE_OFN1584_n_16657
FE_OFN1585_n_16657
FE_OFN1586_n_16657
FE_OFN1587_n_4669
FE_OFN1588_n_4669
FE_OFN1589_n_4669
FE_OFN1590_n_4669
FE_OFN1591_n_4669
FE_OFN1592_n_4669
FE_OFN1593_n_9528
FE_OFN1594_n_9528
FE_OFN1595_n_9528
FE_OFN1596_n_9528
FE_OFN1597_n_9528
FE_OFN1598_n_9528
FE_OFN1599_n_9528
FE_OFN1600_n_9528
FE_OFN1601_n_9528
FE_OFN1602_n_9528
FE_OFN1603_n_9528
FE_OFN1604_n_4740
FE_OFN1607_n_4740
FE_OFN1608_n_4740
FE_OFN1609_n_4740
FE_OFN1610_n_4740
FE_OFN1611_n_4740
FE_OFN1612_n_4740
FE_OFN1613_n_4740
FE_OFN1614_n_4740
FE_OFN1615_n_4740
FE_OFN1616_n_3368
FE_OFN1617_n_3368
FE_OFN1618_n_3368
FE_OFN1620_n_9836
FE_OFN1621_n_9836
FE_OFN1622_n_9836
FE_OFN1623_n_9880
FE_OFN1624_n_9880
FE_OFN1625_n_9880
FE_OFN1626_n_9849
FE_OFN1627_n_9849
FE_OFN1628_n_9849
FE_OFN1629_n_9862
FE_OFN1630_n_9862
FE_OFN1631_n_9862
FE_OFN1632_n_9862
FE_OFN1633_n_16497
FE_OFN1634_n_16497
FE_OFN1635_n_16497
FE_OFN1636_n_16497
FE_OFN1637_n_16497
FE_OFN1638_n_16760
FE_OFN1639_n_16760
FE_OFN1640_n_16760
FE_OFN1641_n_16760
FE_OFN1642_n_16760
FE_OFN1643_n_5751
FE_OFN1644_n_5751
FE_OFN1645_n_5751
FE_OFN1646_n_5751
FE_OFN1647_n_5751
FE_OFN1650_n_4868
FE_OFN1651_n_4868
FE_OFN1652_n_4868
FE_OFN1653_n_4868
FE_OFN1654_n_4868
FE_OFN1655_n_4868
FE_OFN1656_n_4868
FE_OFN1657_n_13650
FE_OFN1658_n_13650
FE_OFN1659_n_13651
FE_OFN1660_n_13651
FE_OFN1663_n_13655
FE_OFN1664_n_13655
FE_OFN1667_n_13664
FE_OFN1668_n_13664
FE_OFN1669_n_13669
FE_OFN1670_n_13669
FE_OFN1671_n_13672
FE_OFN1672_n_13672
FE_OFN1673_n_13673
FE_OFN1674_n_13673
FE_OFN1675_n_10588
FE_OFN1676_n_10588
FE_OFN1677_n_10588
FE_OFN1678_n_10588
FE_OFN1679_n_10588
FE_OFN1680_n_10588
FE_OFN1681_n_16891
FE_OFN1682_n_16891
FE_OFN1683_n_16891
FE_OFN1684_n_16891
FE_OFN1685_n_16891
FE_OFN1686_n_15534
FE_OFN1687_n_15534
FE_OFN1688_n_15534
FE_OFN1689_n_15534
FE_OFN1690_n_15534
FE_OFN1691_n_16992
FE_OFN1692_n_16992
FE_OFN1693_n_16992
FE_OFN1694_n_16992
FE_OFN1695_n_16992
FE_OFN1697_n_9975
FE_OFN1698_n_9975
FE_OFN1699_n_9975
FE_OFN1700_n_9975
FE_OFN1701_n_10892
FE_OFN1702_n_10892
FE_OFN1703_n_10892
FE_OFN1704_n_10892
FE_OFN1705_n_10892
FE_OFN1706_n_10892
FE_OFN1707_n_9320
FE_OFN1708_n_9320
FE_OFN1709_n_9320
FE_OFN1710_n_9320
FE_OFN1712_n_9320
FE_OFN1713_n_9320
FE_OFN1714_n_16637
FE_OFN1715_n_16637
FE_OFN1716_n_16637
FE_OFN1717_n_16637
FE_OFN1718_n_16317
FE_OFN1719_n_16317
FE_OFN1720_n_16317
FE_OFN1722_n_16317
FE_OFN1723_n_16317
FE_OFN1725_n_14987
FE_OFN1726_n_14987
FE_OFN1729_n_11019
FE_OFN1731_n_11019
FE_OFN1732_n_11019
FE_OFN1733_n_11019
FE_OFN1734_n_12004
FE_OFN1736_n_12004
FE_OFN1737_n_12004
FE_OFN1738_n_12004
FE_OFN1739_n_12004
FE_OFN1740_n_12004
FE_OFN1741_n_12086
FE_OFN1743_n_12086
FE_OFN1744_n_12086
FE_OFN1745_n_12086
FE_OFN1746_n_11027
FE_OFN1747_n_11027
FE_OFN1750_n_11027
FE_OFN1751_n_11027
FE_OFN1753_n_12681
FE_OFN1754_n_12681
FE_OFN1755_n_12681
FE_OFN1756_n_13997
FE_OFN1757_n_13997
FE_OFN1759_n_13997
FE_OFN1761_n_14054
FE_OFN1762_n_14054
FE_OFN1763_n_14054
FE_OFN1764_n_14054
FE_OFN1765_n_14054
FE_OFN1766_n_13800
FE_OFN1767_n_13800
FE_OFN1768_n_13800
FE_OFN1770_n_13800
FE_OFN1771_n_13800
FE_OFN1772_n_13800
FE_OFN1773_n_13800
FE_OFN1774_n_13971
FE_OFN1776_n_13971
FE_OFN1777_n_13971
FE_OFN1778_n_13971
FE_OFN1779_wishbone_slave_unit_pci_initiator_if_data_source
FE_OFN1780_wishbone_slave_unit_pci_initiator_if_data_source
FE_OFN1781_wishbone_slave_unit_pci_initiator_if_data_source
FE_OFN1783_wishbone_slave_unit_pci_initiator_if_data_source
FE_OFN1784_wishbone_slave_unit_pci_initiator_if_data_source
FE_OFN1785_wishbone_slave_unit_pci_initiator_if_data_source
FE_OFN1787_n_1699
FE_OFN1788_n_1699
FE_OFN1789_n_1699
FE_OFN1790_n_1699
FE_OFN1791_n_1699
FE_OFN1793_n_4508
FE_OFN1794_n_4508
FE_OFN1795_n_4508
FE_OFN1796_n_4508
FE_OFN1797_n_4508
FE_OFN1798_n_1699
FE_OFN1799_n_1699
FE_OFN179_n_7210
FE_OFN1800_n_1699
FE_OFN1801_n_1699
FE_OFN1803_n_3741
FE_OFN1804_n_3741
FE_OFN1805_n_9899
FE_OFN1806_n_9899
FE_OFN1807_n_9899
FE_OFN1808_n_2047
FE_OFN1809_n_2047
FE_OFN1810_n_2047
FE_OFN1811_n_2047
FE_OFN1812_n_9841
FE_OFN1813_n_9841
FE_OFN1814_n_9839
FE_OFN1815_n_9839
FE_OFN1816_n_9825
FE_OFN1817_n_9825
FE_OFN1818_n_9690
FE_OFN1819_n_9690
FE_OFN181_n_7400
FE_OFN1820_n_9690
FE_OFN1821_n_9690
FE_OFN1822_n_9690
FE_OFN1823_n_9690
FE_OFN1824_n_4490
FE_OFN1825_n_4490
FE_OFN1826_n_4490
FE_OFN1827_n_4454
FE_OFN1828_n_4454
FE_OFN1829_n_4454
FE_OFN1830_n_4454
FE_OFN1831_n_4454
FE_OFN1832_n_2053
FE_OFN1833_n_2053
FE_OFN1834_n_2053
FE_OFN1837_n_2678
FE_OFN1838_n_2678
FE_OFN1839_n_2678
FE_OFN1840_n_9828
FE_OFN1841_n_9828
FE_OFN1842_n_9828
FE_OFN1843_n_8934
FE_OFN1844_n_8934
FE_OFN1845_n_9860
FE_OFN1846_n_9860
FE_OFN1847_n_9860
FE_OFN189_n_1193
FE_OFN193_n_2683
FE_OFN197_n_9230
FE_OFN198_n_9228
FE_OFN199_n_9228
FE_OFN2012_n_13447
FE_OFN2013_n_13447
FE_OFN2014_n_15261
FE_OFN2015_n_15261
FE_OFN2016_n_2520
FE_OFN2017_n_2520
FE_OFN2018_n_3046
FE_OFN2019_n_3046
FE_OFN201_n_9140
FE_OFN202_n_9865
FE_OFN203_n_9865
FE_OFN204_n_9126
FE_OFN205_n_9126
FE_OFN206_n_9858
FE_OFN207_n_9858
FE_OFN208_n_9858
FE_OFN210_n_9858
FE_OFN211_n_9124
FE_OFN212_n_9124
FE_OFN213_n_9856
FE_OFN214_n_9856
FE_OFN215_n_9889
FE_OFN216_n_9889
FE_OFN217_n_9853
FE_OFN218_n_9853
FE_OFN219_n_9846
FE_OFN220_n_9846
FE_OFN222_n_9844
FE_OFN223_n_9122
FE_OFN224_n_9122
FE_OFN225_n_9841
FE_OFN226_n_9841
FE_OFN227_n_9120
FE_OFN228_n_9120
FE_OFN229_n_9839
FE_OFN230_n_9839
FE_OFN231_n_9876
FE_OFN232_n_9876
FE_OFN233_n_9876
FE_OFN234_n_9834
FE_OFN235_n_9834
FE_OFN236_n_9834
FE_OFN237_n_9118
FE_OFN238_n_9118
FE_OFN239_n_9118
FE_OFN240_n_9832
FE_OFN241_n_9832
FE_OFN242_n_9832
FE_OFN243_n_9830
FE_OFN244_n_9830
FE_OFN246_n_9116
FE_OFN248_n_9114
FE_OFN249_n_9112
FE_OFN250_n_9112
FE_OFN251_n_9789
FE_OFN252_n_9789
FE_OFN253_n_9868
FE_OFN254_n_9868
FE_OFN255_n_9825
FE_OFN256_n_9825
FE_OFN257_n_8969
FE_OFN258_n_8969
FE_OFN263_n_9851
FE_OFN264_n_9851
FE_OFN267_n_9884
FE_OFN268_n_9884
FE_OFN273_n_9828
FE_OFN274_n_9828
FE_OFN277_n_9941
FE_OFN278_n_9941
FE_OFN279_n_9941
FE_OFN2_n_4778
FE_OFN319_g66077_p
FE_OFN321_g66081_p
FE_OFN322_g66081_p
FE_OFN323_g66089_p
FE_OFN324_g66089_p
FE_OFN325_g66125_p
FE_OFN416_n_10595
FE_OFN448_n_10853
FE_OFN452_n_10892
FE_OFN487_n_13221
FE_OFN490_n_15978
FE_OFN491_n_15978
FE_OFN492_n_15978
FE_OFN493_n_15978
FE_OFN495_n_9697
FE_OFN496_n_9697
FE_OFN497_n_9697
FE_OFN498_n_9697
FE_OFN499_n_9697
FE_OFN501_n_9697
FE_OFN503_n_9428
FE_OFN505_n_9428
FE_OFN506_n_9899
FE_OFN507_n_9899
FE_OFN508_n_9899
FE_OFN509_n_9899
FE_OFN510_n_9899
FE_OFN511_n_9899
FE_OFN512_n_9899
FE_OFN513_n_9823
FE_OFN514_n_9823
FE_OFN515_n_9823
FE_OFN516_n_9823
FE_OFN517_n_9823
FE_OFN519_n_9690
FE_OFN520_n_9690
FE_OFN521_n_9690
FE_OFN522_n_9690
FE_OFN523_n_9690
FE_OFN524_n_9690
FE_OFN531_n_9864
FE_OFN533_n_9864
FE_OFN534_n_9864
FE_OFN535_n_9895
FE_OFN536_n_9895
FE_OFN537_n_9895
FE_OFN538_n_9895
FE_OFN539_n_9895
FE_OFN540_n_9895
FE_OFN548_n_9502
FE_OFN549_n_9902
FE_OFN550_n_9902
FE_OFN551_n_9902
FE_OFN552_n_9902
FE_OFN554_n_9902
FE_OFN555_n_9902
FE_OFN557_n_9531
FE_OFN559_n_9531
FE_OFN560_n_9531
FE_OFN561_n_9692
FE_OFN562_n_9692
FE_OFN563_n_9692
FE_OFN564_n_9692
FE_OFN565_n_9692
FE_OFN566_n_9692
FE_OFN567_n_9694
FE_OFN568_n_9694
FE_OFN569_n_9694
FE_OFN570_n_9694
FE_OFN571_n_9694
FE_OFN572_n_9694
FE_OFN573_n_9687
FE_OFN574_n_9687
FE_OFN575_n_9687
FE_OFN576_n_9687
FE_OFN577_n_9687
FE_OFN579_n_9904
FE_OFN580_n_9904
FE_OFN581_n_9904
FE_OFN588_n_4490
FE_OFN589_n_4490
FE_OFN590_n_4490
FE_OFN591_n_4490
FE_OFN593_n_4409
FE_OFN594_n_4409
FE_OFN595_n_4409
FE_OFN596_n_4409
FE_OFN597_n_4409
FE_OFN598_n_4454
FE_OFN599_n_4454
FE_OFN600_n_4454
FE_OFN601_n_4454
FE_OFN602_n_4454
FE_OFN605_n_4669
FE_OFN607_n_4669
FE_OFN611_n_4497
FE_OFN612_n_4497
FE_OFN613_n_4497
FE_OFN614_n_4497
FE_OFN615_n_4497
FE_OFN621_n_4671
FE_OFN624_n_4392
FE_OFN625_n_4392
FE_OFN626_n_4392
FE_OFN627_n_4392
FE_OFN628_n_4495
FE_OFN629_n_4495
FE_OFN630_n_4495
FE_OFN631_n_4495
FE_OFN632_n_4495
FE_OFN633_n_4505
FE_OFN634_n_4505
FE_OFN635_n_4505
FE_OFN636_n_4505
FE_OFN637_n_4505
FE_OFN640_n_4655
FE_OFN644_n_4460
FE_OFN647_n_4460
FE_OFN649_n_4417
FE_OFN650_n_4417
FE_OFN651_n_4417
FE_OFN652_n_4417
FE_OFN653_n_4417
FE_OFN654_n_4438
FE_OFN655_n_4438
FE_OFN656_n_4438
FE_OFN657_n_4438
FE_OFN658_n_4438
FE_OFN667_n_8232
FE_OFN668_n_8232
FE_OFN669_n_8232
FE_OFN670_n_8232
FE_OFN671_n_8232
FE_OFN672_n_8232
FE_OFN673_n_8140
FE_OFN674_n_8140
FE_OFN675_n_8140
FE_OFN678_n_8060
FE_OFN679_n_8060
FE_OFN680_n_8060
FE_OFN688_n_7350
FE_OFN698_n_7498
FE_OFN709_n_16779
FE_OFN716_n_11795
FE_OFN717_n_11795
FE_OFN719_n_11138
FE_OFN723_n_9163
FE_OFN724_n_9163
FE_OFN734_n_15366
FE_OFN735_n_15366
FE_OFN736_n_15366
FE_OFN737_n_4152
FE_OFN738_n_4152
FE_OFN741_n_2678
FE_OFN743_n_2678
FE_OFN747_n_2678
FE_OFN748_n_2678
FE_OFN751_n_2547
FE_OFN752_n_2547
FE_OFN753_n_2520
FE_OFN754_n_2520
FE_OFN7_n_11877
FE_OFN852_n_4736
FE_OFN853_n_4736
FE_OFN854_n_4736
FE_OFN855_n_4736
FE_OFN856_n_4734
FE_OFN857_n_4734
FE_OFN858_n_4734
FE_OFN859_n_4734
FE_OFN860_n_4734
FE_OFN868_n_4725
FE_OFN869_n_4725
FE_OFN887_n_2292
FE_OFN888_n_2292
FE_OFN889_n_2292
FE_OFN890_n_2292
FE_OFN891_n_2292
FE_OFN892_n_2047
FE_OFN893_n_2047
FE_OFN894_n_2047
FE_OFN895_n_2047
FE_OFN896_n_2047
FE_OFN897_n_2248
FE_OFN898_n_2248
FE_OFN899_n_2248
FE_OFN8_n_11877
FE_OFN900_n_2248
FE_OFN901_n_2055
FE_OFN902_n_2055
FE_OFN903_n_2055
FE_OFN904_n_2055
FE_OFN906_n_1699
FE_OFN907_n_1699
FE_OFN909_n_2299
FE_OFN910_n_2299
FE_OFN911_n_2299
FE_OFN912_n_2299
FE_OFN913_n_2053
FE_OFN914_n_2053
FE_OFN916_n_2053
FE_OFN924_n_13784
FE_OFN931_n_2700
FE_OFN933_n_2697
FE_OFN934_n_2697
FE_OFN935_n_2696
FE_OFN937_n_574
FE_OFN938_n_574
FE_OFN939_n_574
FE_OFN940_n_16089
FE_OFN941_n_16089
FE_OFN942_n_16288
FE_OFN943_n_16288
FE_OFN944_n_16288
FE_OFN945_n_16288
FE_OFN946_n_16288
FE_OFN949_n_4725
FE_OFN950_n_4725
FE_OFN951_n_4725
FE_OFN952_n_4725
FE_OFN953_n_4725
FE_OFN954_n_1036
FE_OFN956_n_11877
FE_OFN959_n_16760
FE_OFN962_n_16810
FE_OFN965_n_4655
FE_OFN966_n_4655
FE_OFN967_n_4655
FE_OFN968_n_4655
FE_OFN969_n_4655
FE_OFN970_n_4727
FE_OFN973_n_4727
FE_OFN974_n_4727
FE_OFN975_n_4727
FE_OFN976_n_4727
FE_OFN977_n_4727
FE_OFN978_n_4727
FE_OFN979_n_7102
FE_OFN980_n_7102
FE_OFN981_n_7102
FE_OFN984_n_16720
FE_OFN986_n_16720
FE_OFN987_n_15729
FE_OFN988_n_15729
FE_OFN989_n_15729
FE_OFN990_n_15729
FE_OFN991_n_15729
FE_OFN993_n_4778
FE_OFN994_n_4778
FE_OFN995_n_4778
FE_OFN996_n_7350
FE_OFN997_n_7350
FE_OFN998_n_7350
FE_OFN999_n_7350
FE_OFN99_n_12086
FE_RN_0_0
FE_RN_102_0
FE_RN_103_0
FE_RN_104_0
FE_RN_105_0
FE_RN_106_0
FE_RN_107_0
FE_RN_108_0
FE_RN_109_0
FE_RN_110_0
FE_RN_111_0
FE_RN_112_0
FE_RN_113_0
FE_RN_114_0
FE_RN_115_0
FE_RN_116_0
FE_RN_117_0
FE_RN_118_0
FE_RN_119_0
FE_RN_11_0
FE_RN_120_0
FE_RN_121_0
FE_RN_122_0
FE_RN_123_0
FE_RN_126_0
FE_RN_127_0
FE_RN_128_0
FE_RN_129_0
FE_RN_130_0
FE_RN_131_0
FE_RN_132_0
FE_RN_133_0
FE_RN_134_0
FE_RN_137_0
FE_RN_138_0
FE_RN_139_0
FE_RN_140_0
FE_RN_141_0
FE_RN_142_0
FE_RN_143_0
FE_RN_150_0
FE_RN_151_0
FE_RN_152_0
FE_RN_156_0
FE_RN_157_0
FE_RN_158_0
FE_RN_159_0
FE_RN_15_0
FE_RN_160_0
FE_RN_161_0
FE_RN_162_0
FE_RN_163_0
FE_RN_164_0
FE_RN_171_0
FE_RN_172_0
FE_RN_173_0
FE_RN_174_0
FE_RN_175_0
FE_RN_176_0
FE_RN_177_0
FE_RN_178_0
FE_RN_179_0
FE_RN_17_0
FE_RN_180_0
FE_RN_182_0
FE_RN_188_0
FE_RN_189_0
FE_RN_190_0
FE_RN_191_0
FE_RN_192_0
FE_RN_193_0
FE_RN_194_0
FE_RN_198_0
FE_RN_199_0
FE_RN_1_0
FE_RN_200_0
FE_RN_201_0
FE_RN_202_0
FE_RN_203_0
FE_RN_204_0
FE_RN_205_0
FE_RN_206_0
FE_RN_207_0
FE_RN_208_0
FE_RN_209_0
FE_RN_213_0
FE_RN_214_0
FE_RN_215_0
FE_RN_216_0
FE_RN_217_0
FE_RN_218_0
FE_RN_219_0
FE_RN_220_0
FE_RN_221_0
FE_RN_222_0
FE_RN_223_0
FE_RN_224_0
FE_RN_226_0
FE_RN_227_0
FE_RN_228_0
FE_RN_229_0
FE_RN_230_0
FE_RN_231_0
FE_RN_232_0
FE_RN_233_0
FE_RN_234_0
FE_RN_239_0
FE_RN_241_0
FE_RN_242_0
FE_RN_243_0
FE_RN_245_0
FE_RN_24_0
FE_RN_251_0
FE_RN_252_0
FE_RN_253_0
FE_RN_254_0
FE_RN_255_0
FE_RN_256_0
FE_RN_257_0
FE_RN_258_0
FE_RN_25_0
FE_RN_260_0
FE_RN_261_0
FE_RN_262_0
FE_RN_263_0
FE_RN_264_0
FE_RN_265_0
FE_RN_266_0
FE_RN_267_0
FE_RN_268_0
FE_RN_269_0
FE_RN_26_0
FE_RN_270_0
FE_RN_271_0
FE_RN_272_0
FE_RN_273_0
FE_RN_274_0
FE_RN_283_0
FE_RN_284_0
FE_RN_285_0
FE_RN_286_0
FE_RN_292_0
FE_RN_293_0
FE_RN_294_0
FE_RN_297_0
FE_RN_298_0
FE_RN_299_0
FE_RN_2_0
FE_RN_300_0
FE_RN_301_0
FE_RN_302_0
FE_RN_307_0
FE_RN_308_0
FE_RN_309_0
FE_RN_30_0
FE_RN_310_0
FE_RN_311_0
FE_RN_312_0
FE_RN_313_0
FE_RN_315_0
FE_RN_316_0
FE_RN_318_0
FE_RN_31_0
FE_RN_323_0
FE_RN_324_0
FE_RN_325_0
FE_RN_326_0
FE_RN_327_0
FE_RN_328_0
FE_RN_32_0
FE_RN_331_0
FE_RN_332_0
FE_RN_333_0
FE_RN_334_0
FE_RN_335_0
FE_RN_336_0
FE_RN_337_0
FE_RN_338_0
FE_RN_339_0
FE_RN_33_0
FE_RN_340_0
FE_RN_341_0
FE_RN_342_0
FE_RN_344_0
FE_RN_345_0
FE_RN_34_0
FE_RN_350_0
FE_RN_351_0
FE_RN_352_0
FE_RN_353_0
FE_RN_354_0
FE_RN_355_0
FE_RN_356_0
FE_RN_358_0
FE_RN_359_0
FE_RN_35_0
FE_RN_360_0
FE_RN_361_0
FE_RN_362_0
FE_RN_363_0
FE_RN_364_0
FE_RN_369_0
FE_RN_36_0
FE_RN_371_0
FE_RN_372_0
FE_RN_373_0
FE_RN_377_0
FE_RN_378_0
FE_RN_37_0
FE_RN_381_0
FE_RN_38_0
FE_RN_391_0
FE_RN_392_0
FE_RN_393_0
FE_RN_394_0
FE_RN_395_0
FE_RN_396_0
FE_RN_399_0
FE_RN_39_0
FE_RN_3_0
FE_RN_402_0
FE_RN_403_0
FE_RN_404_0
FE_RN_405_0
FE_RN_40_0
FE_RN_41_0
FE_RN_427_0
FE_RN_42_0
FE_RN_430_0
FE_RN_431_0
FE_RN_432_0
FE_RN_433_0
FE_RN_434_0
FE_RN_435_0
FE_RN_436_0
FE_RN_437_0
FE_RN_438_0
FE_RN_439_0
FE_RN_43_0
FE_RN_440_0
FE_RN_441_0
FE_RN_442_0
FE_RN_443_0
FE_RN_444_0
FE_RN_445_0
FE_RN_446_0
FE_RN_447_0
FE_RN_448_0
FE_RN_449_0
FE_RN_44_0
FE_RN_451_0
FE_RN_45_0
FE_RN_46_0
FE_RN_47_0
FE_RN_48_0
FE_RN_49_0
FE_RN_4_0
FE_RN_50_0
FE_RN_51_0
FE_RN_52_0
FE_RN_53_0
FE_RN_58_0
FE_RN_59_0
FE_RN_5_0
FE_RN_60_0
FE_RN_61_0
FE_RN_62_0
FE_RN_63_0
FE_RN_64_0
FE_RN_65_0
FE_RN_66_0
FE_RN_67_0
FE_RN_68_0
FE_RN_69_0
FE_RN_70_0
FE_RN_71_0
FE_RN_72_0
FE_RN_73_0
FE_RN_74_0
FE_RN_75_0
FE_RN_76_0
FE_RN_77_0
FE_RN_78_0
FE_RN_79_0
FE_RN_80_0
FE_RN_81_0
FE_RN_82_0
FE_RN_83_0
FE_RN_85_0
FE_RN_87_0
FE_RN_88_0
FE_RN_89_0
FE_RN_90_0
FE_RN_91_0
FE_RN_92_0
FE_RN_96_0
FE_RN_97_0
FE_RN_98_0
FE_RN_99_0
FE_RN_9_0
conf_pci_init_complete_out
conf_target_abort_recv_in
conf_w_addr_in
conf_w_addr_in_931
conf_w_addr_in_932
conf_w_addr_in_933
conf_w_addr_in_935
conf_w_addr_in_937
conf_w_addr_in_938
conf_w_addr_in_939
conf_wb_err_addr_in_943
conf_wb_err_addr_in_944
conf_wb_err_addr_in_945
conf_wb_err_addr_in_946
conf_wb_err_addr_in_947
conf_wb_err_addr_in_948
conf_wb_err_addr_in_949
conf_wb_err_addr_in_950
conf_wb_err_addr_in_951
conf_wb_err_addr_in_952
conf_wb_err_addr_in_953
conf_wb_err_addr_in_954
conf_wb_err_addr_in_955
conf_wb_err_addr_in_956
conf_wb_err_addr_in_957
conf_wb_err_addr_in_958
conf_wb_err_addr_in_959
conf_wb_err_addr_in_960
conf_wb_err_addr_in_961
conf_wb_err_addr_in_962
conf_wb_err_addr_in_963
conf_wb_err_addr_in_964
conf_wb_err_addr_in_965
conf_wb_err_addr_in_966
conf_wb_err_addr_in_967
conf_wb_err_addr_in_968
conf_wb_err_addr_in_969
conf_wb_err_addr_in_970
conf_wb_err_addr_in_971
conf_wb_err_bc_in
conf_wb_err_bc_in_848
configuration_cache_line_size_reg
configuration_cache_line_size_reg_2996
configuration_int_meta
configuration_interrupt_line
configuration_interrupt_line_37
configuration_interrupt_line_38
configuration_interrupt_line_39
configuration_interrupt_line_40
configuration_interrupt_line_41
configuration_interrupt_line_42
configuration_interrupt_line_43
configuration_interrupt_out_reg_Q
configuration_meta_cache_lsize_to_wb_bits
configuration_meta_cache_lsize_to_wb_bits_926
configuration_meta_cache_lsize_to_wb_bits_930
configuration_meta_cache_lsize_to_wb_bits_931
configuration_meta_pci_err_cs_bits
configuration_pci_err_addr_471
configuration_pci_err_addr_472
configuration_pci_err_addr_473
configuration_pci_err_addr_475
configuration_pci_err_addr_476
configuration_pci_err_addr_477
configuration_pci_err_addr_478
configuration_pci_err_addr_481
configuration_pci_err_addr_482
configuration_pci_err_addr_483
configuration_pci_err_addr_484
configuration_pci_err_addr_485
configuration_pci_err_addr_486
configuration_pci_err_addr_487
configuration_pci_err_addr_488
configuration_pci_err_addr_489
configuration_pci_err_addr_490
configuration_pci_err_addr_491
configuration_pci_err_addr_492
configuration_pci_err_addr_493
configuration_pci_err_addr_494
configuration_pci_err_addr_495
configuration_pci_err_addr_496
configuration_pci_err_addr_497
configuration_pci_err_addr_498
configuration_pci_err_addr_499
configuration_pci_err_addr_500
configuration_pci_err_addr_501
configuration_pci_err_cs_bit0
configuration_pci_err_cs_bit10
configuration_pci_err_cs_bit31_24
configuration_pci_err_cs_bit8
configuration_pci_err_cs_bit9
configuration_pci_err_cs_bit_464
configuration_pci_err_cs_bit_465
configuration_pci_err_cs_bit_466
configuration_pci_err_cs_bit_467
configuration_pci_err_cs_bit_468
configuration_pci_err_cs_bit_469
configuration_pci_err_cs_bit_470
configuration_pci_err_data
configuration_pci_err_data_502
configuration_pci_err_data_503
configuration_pci_err_data_504
configuration_pci_err_data_506
configuration_pci_err_data_508
configuration_pci_err_data_510
configuration_pci_err_data_511
configuration_pci_err_data_513
configuration_pci_err_data_514
configuration_pci_err_data_515
configuration_pci_err_data_516
configuration_pci_err_data_517
configuration_pci_err_data_518
configuration_pci_err_data_519
configuration_pci_err_data_520
configuration_pci_err_data_521
configuration_pci_err_data_522
configuration_pci_err_data_524
configuration_pci_err_data_525
configuration_pci_err_data_526
configuration_pci_err_data_527
configuration_pci_err_data_528
configuration_pci_err_data_529
configuration_pci_err_data_530
configuration_pci_err_data_531
configuration_pci_err_data_532
configuration_rst_inactive
configuration_rst_inactive_sync
configuration_set_pci_err_cs_bit8
configuration_set_pci_err_cs_bit8_reg_Q
configuration_status_bit8
configuration_status_bit_322
configuration_status_bit_351
configuration_status_bit_379
configuration_status_bit_407
configuration_status_bit_435
configuration_sync_cache_lsize_to_wb_bits_reg_2__Q
configuration_sync_cache_lsize_to_wb_bits_reg_3__Q
configuration_sync_command_bit0
configuration_sync_command_bit1
configuration_sync_command_bit2
configuration_sync_command_bit6
configuration_sync_command_bit8
configuration_sync_init_complete
configuration_sync_pci_err_cs_8_del_bit_reg_Q
configuration_sync_pci_err_cs_8_delayed_bckp_bit
configuration_sync_pci_err_cs_8_delayed_bckp_bit_reg_Q
configuration_sync_pci_err_cs_8_meta_bckp_bit
configuration_sync_pci_err_cs_8_meta_del_bit
configuration_sync_pci_err_cs_8_sync_bckp_bit
configuration_wb_err_addr_533
configuration_wb_err_addr_534
configuration_wb_err_addr_535
configuration_wb_err_addr_536
configuration_wb_err_addr_537
configuration_wb_err_addr_538
configuration_wb_err_addr_540
configuration_wb_err_addr_541
configuration_wb_err_addr_542
configuration_wb_err_addr_543
configuration_wb_err_addr_544
configuration_wb_err_addr_545
configuration_wb_err_addr_546
configuration_wb_err_addr_547
configuration_wb_err_addr_548
configuration_wb_err_addr_549
configuration_wb_err_addr_550
configuration_wb_err_addr_551
configuration_wb_err_addr_552
configuration_wb_err_addr_553
configuration_wb_err_addr_554
configuration_wb_err_addr_555
configuration_wb_err_addr_556
configuration_wb_err_addr_558
configuration_wb_err_addr_559
configuration_wb_err_addr_560
configuration_wb_err_addr_561
configuration_wb_err_addr_562
configuration_wb_err_addr_563
configuration_wb_err_cs_bit0
configuration_wb_err_cs_bit31_24
configuration_wb_err_cs_bit_564
configuration_wb_err_cs_bit_565
configuration_wb_err_cs_bit_566
configuration_wb_err_cs_bit_567
configuration_wb_err_cs_bit_568
configuration_wb_err_cs_bit_569
configuration_wb_err_cs_bit_570
configuration_wb_err_data
configuration_wb_err_data_572
configuration_wb_err_data_573
configuration_wb_err_data_574
configuration_wb_err_data_578
configuration_wb_err_data_579
configuration_wb_err_data_581
configuration_wb_err_data_582
configuration_wb_err_data_583
configuration_wb_err_data_584
configuration_wb_err_data_585
configuration_wb_err_data_586
configuration_wb_err_data_587
configuration_wb_err_data_588
configuration_wb_err_data_589
configuration_wb_err_data_590
configuration_wb_err_data_591
configuration_wb_err_data_592
configuration_wb_err_data_593
configuration_wb_err_data_594
configuration_wb_err_data_595
configuration_wb_err_data_596
configuration_wb_err_data_597
configuration_wb_err_data_598
configuration_wb_err_data_599
configuration_wb_err_data_600
configuration_wb_err_data_601
g20_dup74712_db
g22_p
g52252_p
g52253_p
g52393_da
g52393_db
g52393_sb
g52394_da
g52394_db
g52394_sb
g52395_da
g52395_db
g52395_sb
g52396_da
g52396_db
g52396_sb
g52397_da
g52397_db
g52397_sb
g52398_da
g52398_db
g52398_sb
g52399_da
g52399_db
g52399_sb
g52400_da
g52400_db
g52400_sb
g52401_da
g52401_db
g52401_sb
g52402_da
g52402_db
g52402_sb
g52403_da
g52403_db
g52403_sb
g52404_da
g52404_db
g52404_sb
g52405_da
g52405_db
g52405_sb
g52439_da
g52439_db
g52440_da
g52440_db
g52440_sb
g52441_da
g52441_db
g52441_sb
g52442_da
g52442_db
g52442_sb
g52443_da
g52443_db
g52443_sb
g52444_da
g52444_db
g52444_sb
g52445_da
g52445_db
g52446_da
g52446_db
g52446_sb
g52447_da
g52447_db
g52447_sb
g52448_da
g52448_db
g52448_sb
g52449_da
g52449_db
g52449_sb
g52450_da
g52450_db
g52450_sb
g52451_da
g52451_db
g52451_sb
g52452_da
g52452_db
g52452_sb
g52453_da
g52453_db
g52453_sb
g52454_da
g52454_db
g52454_sb
g52455_da
g52455_db
g52455_sb
g52456_da
g52456_db
g52456_sb
g52457_da
g52457_db
g52457_sb
g52458_da
g52458_db
g52458_sb
g52459_da
g52459_db
g52459_sb
g52460_da
g52460_db
g52460_sb
g52461_da
g52461_db
g52461_sb
g52462_da
g52462_db
g52462_sb
g52463_da
g52463_db
g52463_sb
g52464_da
g52464_db
g52464_sb
g52465_da
g52465_db
g52465_sb
g52466_da
g52466_db
g52466_sb
g52467_da
g52467_db
g52467_sb
g52468_da
g52468_db
g52468_sb
g52469_da
g52469_db
g52469_sb
g52470_da
g52470_db
g52470_sb
g52471_da
g52471_db
g52471_sb
g52472_da
g52472_db
g52472_sb
g52473_da
g52473_db
g52473_sb
g52474_da
g52474_db
g52474_sb
g52475_da
g52475_db
g52475_sb
g52476_da
g52476_db
g52476_sb
g52477_da
g52477_db
g52477_sb
g52478_da
g52478_db
g52478_sb
g52479_da
g52479_db
g52480_da
g52480_db
g52480_sb
g52481_da
g52481_db
g52482_da
g52482_db
g52482_sb
g52483_da
g52483_db
g52483_sb
g52484_da
g52484_sb
g52485_da
g52485_db
g52485_sb
g52495_p
g52496_p
g52497_p
g52498_p
g52503_da
g52503_db
g52503_sb
g52504_da
g52504_db
g52504_sb
g52505_da
g52505_db
g52505_sb
g52506_da
g52506_db
g52506_sb
g52507_da
g52507_db
g52507_sb
g52508_da
g52508_db
g52508_sb
g52509_da
g52509_db
g52509_sb
g52510_da
g52510_db
g52510_sb
g52511_da
g52511_db
g52511_sb
g52512_da
g52512_db
g52512_sb
g52513_da
g52513_db
g52513_sb
g52514_da
g52514_db
g52514_sb
g52515_da
g52515_db
g52515_sb
g52516_da
g52516_db
g52516_sb
g52517_da
g52517_db
g52517_sb
g52518_da
g52518_db
g52518_sb
g52519_da
g52519_db
g52519_sb
g52520_da
g52520_db
g52520_sb
g52521_da
g52521_db
g52521_sb
g52522_da
g52522_db
g52522_sb
g52523_da
g52523_db
g52523_sb
g52524_da
g52524_db
g52524_sb
g52525_da
g52525_db
g52525_sb
g52526_da
g52526_db
g52526_sb
g52527_da
g52527_db
g52527_sb
g52529_da
g52529_db
g52529_sb
g52530_da
g52530_db
g52530_sb
g52531_da
g52531_db
g52531_sb
g52532_da
g52532_db
g52532_sb
g52533_da
g52533_db
g52533_sb
g52534_da
g52534_db
g52534_sb
g52590_da
g52590_db
g52590_sb
g52591_da
g52591_db
g52591_sb
g52592_da
g52592_db
g52592_sb
g52593_da
g52593_db
g52593_sb
g52594_da
g52594_db
g52594_sb
g52595_da
g52595_db
g52595_sb
g52596_da
g52596_db
g52596_sb
g52597_da
g52597_db
g52597_sb
g52598_da
g52598_db
g52598_sb
g52599_da
g52599_db
g52599_sb
g52600_da
g52600_db
g52600_sb
g52601_da
g52601_db
g52601_sb
g52602_da
g52602_db
g52602_sb
g52603_da
g52603_db
g52603_sb
g52604_da
g52604_db
g52604_sb
g52605_da
g52605_db
g52605_sb
g52606_da
g52606_db
g52606_sb
g52607_da
g52607_db
g52607_sb
g52608_da
g52608_db
g52608_sb
g52609_da
g52609_db
g52609_sb
g52610_da
g52610_db
g52610_sb
g52611_da
g52611_db
g52611_sb
g52612_da
g52612_db
g52612_sb
g52614_da
g52614_db
g52614_sb
g52616_da
g52616_db
g52616_sb
g52617_da
g52617_db
g52617_sb
g52618_da
g52618_db
g52618_sb
g52619_da
g52619_db
g52619_sb
g52620_da
g52620_db
g52620_sb
g52621_da
g52621_db
g52621_sb
g52622_da
g52622_db
g52622_sb
g52623_p
g52624_da
g52624_db
g52624_sb
g52625_da
g52625_db
g52625_sb
g52626_da
g52626_db
g52627_da
g52627_db
g52627_sb
g52628_da
g52628_db
g52628_sb
g52629_da
g52629_db
g52629_sb
g52630_da
g52630_db
g52630_sb
g52631_da
g52631_db
g52631_sb
g52632_da
g52632_db
g52632_sb
g52633_da
g52633_db
g52633_sb
g52634_da
g52634_db
g52634_sb
g52635_da
g52635_db
g52635_sb
g52636_da
g52636_db
g52636_sb
g52637_da
g52637_db
g52639_da
g52639_db
g52640_da
g52640_db
g52640_sb
g52641_da
g52641_db
g52641_sb
g52642_da
g52642_db
g52642_sb
g52643_da
g52643_db
g52643_sb
g52644_da
g52644_db
g52644_sb
g52645_da
g52645_db
g52645_sb
g52646_da
g52646_db
g52647_da
g52647_db
g52647_sb
g52648_da
g52648_db
g52648_sb
g52650_da
g52650_db
g52650_sb
g52651_da
g52651_db
g52651_sb
g52652_da
g52652_db
g52653_da
g52653_db
g52653_sb
g52675_p
g52714_p
g52865_p
g52_p
g53011_p
g53012_p
g53014_p
g53017_p
g53018_p
g53022_p
g53026_p
g53031_p
g53035_p
g53039_p
g53069_p
g53071_p
g53072_p
g53073_p
g53074_p
g53076_p
g53077_p
g53078_p
g53079_p
g53080_p
g53082_p
g53083_p
g53105_da
g53105_db
g53105_sb
g53141_p
g53142_p
g53154_p
g53158_p
g53159_p
g53162_p
g53163_p
g53186_p
g53187_p
g53198_p
g53202_p
g53203_p
g53210_p
g53211_p
g53214_p
g53215_p
g53222_p
g53223_p
g53226_p
g53227_p
g53238_p
g53239_p
g53242_p
g53243_p
g53246_p
g53247_p
g53254_p
g53255_p
g53258_p
g53259_p
g53262_p
g53263_p
g53275_p
g53276_p
g53289_p
g53301_p
g53302_p
g53309_p
g53310_p
g53709_p
g53729_p
g53752_p
g53890_da
g53890_db
g53890_sb
g53892_da
g53892_db
g53892_sb
g53897_da
g53897_db
g53897_sb
g53899_da
g53899_db
g53899_sb
g53901_da
g53901_db
g53901_sb
g53902_da
g53902_db
g53902_sb
g53903_da
g53903_db
g53903_sb
g53905_da
g53905_db
g53905_sb
g53906_da
g53906_db
g53906_sb
g53907_da
g53907_db
g53907_sb
g53908_da
g53908_db
g53908_sb
g53909_da
g53909_db
g53909_sb
g53910_da
g53910_db
g53910_sb
g53912_da
g53912_db
g53912_sb
g53913_da
g53913_db
g53913_sb
g53914_da
g53914_db
g53914_sb
g53916_da
g53916_db
g53916_sb
g53918_da
g53918_db
g53918_sb
g53920_da
g53920_db
g53920_sb
g53921_da
g53921_db
g53921_sb
g53922_da
g53922_db
g53922_sb
g53924_da
g53924_db
g53924_sb
g53925_da
g53925_db
g53925_sb
g53926_da
g53926_db
g53926_sb
g53927_da
g53927_sb
g53928_da
g53928_db
g53928_sb
g53929_da
g53929_db
g53929_sb
g53936_da
g53936_db
g53937_da
g53937_db
g53938_da
g53938_db
g53939_da
g53940_da
g53940_db
g53940_sb
g53941_da
g53941_db
g53942_da
g53942_db
g53942_sb
g53943_sb
g53944_da
g53944_db
g53944_sb
g53946_da
g53946_db
g53946_sb
g53947_da
g53947_db
g53990_p
g54030_da
g54030_db
g54030_sb
g54038_db
g54039_da
g54039_db
g54040_da
g54040_db
g54131_da
g54131_sb
g54132_da
g54132_db
g54132_sb
g54133_da
g54133_db
g54133_sb
g54134_da
g54134_db
g54134_sb
g54135_da
g54135_db
g54135_sb
g54137_da
g54137_db
g54137_sb
g54138_da
g54138_db
g54138_sb
g54141_da
g54141_db
g54141_sb
g54142_da
g54142_db
g54143_da
g54143_db
g54145_da
g54145_db
g54145_sb
g54146_da
g54146_db
g54146_sb
g54147_da
g54147_db
g54147_sb
g54149_da
g54149_db
g54149_sb
g54150_da
g54150_db
g54150_sb
g54152_da
g54152_db
g54152_sb
g54153_da
g54153_db
g54153_sb
g54154_da
g54154_db
g54154_sb
g54157_da
g54157_db
g54157_sb
g54161_da
g54161_db
g54161_sb
g54163_da
g54163_db
g54163_sb
g54167_da
g54167_db
g54167_sb
g54169_da
g54169_sb
g54171_da
g54171_db
g54171_sb
g54174_db
g54176_da
g54176_db
g54176_sb
g54177_da
g54177_db
g54177_sb
g54178_da
g54178_db
g54178_sb
g54179_da
g54179_db
g54179_sb
g54180_da
g54180_db
g54180_sb
g54181_da
g54181_db
g54181_sb
g54183_da
g54183_db
g54183_sb
g54185_db
g54186_da
g54186_db
g54186_sb
g54187_da
g54187_db
g54187_sb
g54188_db
g54190_da
g54190_db
g54190_sb
g54191_da
g54191_db
g54191_sb
g54192_da
g54192_db
g54192_sb
g54193_da
g54193_db
g54193_sb
g54194_da
g54194_db
g54194_sb
g54200_da
g54200_db
g54200_sb
g54201_da
g54201_db
g54201_sb
g54202_da
g54202_db
g54202_sb
g54203_da
g54203_db
g54203_sb
g54204_da
g54204_db
g54204_sb
g54205_da
g54205_db
g54205_sb
g54206_da
g54206_db
g54208_da
g54208_db
g54209_da
g54209_db
g54209_sb
g54210_da
g54210_db
g54211_da
g54211_db
g54212_da
g54212_db
g54214_da
g54214_db
g54215_da
g54215_db
g54216_db
g54218_da
g54218_db
g54221_da
g54221_db
g54222_da
g54222_db
g54223_da
g54223_db
g54225_da
g54225_db
g54226_da
g54226_db
g54228_da
g54228_db
g54229_da
g54229_db
g54234_da
g54234_db
g54234_sb
g54235_da
g54235_db
g54235_sb
g54236_da
g54236_db
g54236_sb
g54238_da
g54238_db
g54238_sb
g54239_da
g54239_db
g54239_sb
g54244_db
g54304_da
g54304_db
g54304_sb
g54305_da
g54305_db
g54305_sb
g54306_da
g54306_db
g54306_sb
g54307_da
g54307_db
g54307_sb
g54309_da
g54309_db
g54309_sb
g54310_da
g54310_db
g54310_sb
g54311_da
g54311_db
g54311_sb
g54312_da
g54312_db
g54312_sb
g54313_da
g54313_db
g54313_sb
g54314_da
g54314_db
g54314_sb
g54315_da
g54315_db
g54315_sb
g54316_da
g54316_db
g54316_sb
g54317_da
g54317_db
g54317_sb
g54318_da
g54318_db
g54318_sb
g54319_da
g54319_db
g54319_sb
g54320_da
g54320_db
g54320_sb
g54321_da
g54321_db
g54321_sb
g54322_da
g54322_db
g54322_sb
g54323_da
g54323_db
g54323_sb
g54324_da
g54324_db
g54324_sb
g54325_da
g54325_db
g54325_sb
g54326_da
g54326_db
g54326_sb
g54327_da
g54327_db
g54327_sb
g54328_da
g54328_db
g54328_sb
g54329_p
g54330_da
g54330_db
g54330_sb
g54331_da
g54331_db
g54331_sb
g54332_da
g54332_db
g54332_sb
g54333_da
g54333_db
g54333_sb
g54334_da
g54334_db
g54334_sb
g54335_da
g54335_db
g54335_sb
g54336_da
g54336_db
g54336_sb
g54337_da
g54337_db
g54337_sb
g54338_da
g54338_db
g54338_sb
g54339_da
g54339_db
g54339_sb
g54340_da
g54340_db
g54340_sb
g54341_da
g54341_db
g54341_sb
g54342_da
g54342_db
g54342_sb
g54343_da
g54343_db
g54343_sb
g54344_da
g54344_db
g54344_sb
g54345_da
g54345_db
g54345_sb
g54346_da
g54346_db
g54347_da
g54347_db
g54347_sb
g54348_da
g54348_db
g54348_sb
g54349_da
g54349_db
g54349_sb
g54350_da
g54350_db
g54350_sb
g54351_da
g54351_db
g54351_sb
g54352_da
g54352_db
g54352_sb
g54353_da
g54353_db
g54353_sb
g54354_da
g54354_db
g54354_sb
g54355_da
g54355_db
g54355_sb
g54356_da
g54356_db
g54356_sb
g54357_da
g54357_db
g54357_sb
g54358_da
g54358_db
g54358_sb
g54359_da
g54359_db
g54359_sb
g54360_da
g54360_db
g54360_sb
g54361_da
g54361_db
g54361_sb
g54362_da
g54362_db
g54362_sb
g54363_da
g54363_db
g54363_sb
g54364_da
g54364_db
g54364_sb
g54365_da
g54365_db
g54365_sb
g54366_da
g54366_db
g54366_sb
g54367_da
g54367_db
g54367_sb
g54368_da
g54368_db
g54368_sb
g54369_da
g54369_db
g54369_sb
g54453_p
g54455_p
g54456_p
g54458_p
g54465_p
g54471_da
g54471_db
g54471_sb
g54472_da
g54472_db
g54472_sb
g54484_da
g54484_db
g54484_sb
g54485_da
g54485_db
g54485_sb
g54486_da
g54486_db
g54486_sb
g54487_da
g54487_db
g54487_sb
g54488_da
g54488_db
g54488_sb
g54489_da
g54489_db
g54489_sb
g54490_da
g54490_db
g54490_sb
g54491_da
g54491_db
g54491_sb
g54492_da
g54492_db
g54492_sb
g54493_da
g54493_db
g54493_sb
g54494_da
g54494_db
g54494_sb
g54495_da
g54495_db
g54495_sb
g54572_p
g54573_p
g54574_p
g54579_p
g54580_p
g54581_p
g54587_p
g54593_p
g54595_p
g54597_p
g54601_p
g55851_da
g55851_db
g55851_sb
g55852_da
g55852_db
g55852_sb
g55853_da
g55853_db
g55853_sb
g56933_da
g56933_db
g56933_sb
g56934_da
g56934_db
g56934_sb
g57030_p
g57034_da
g57034_db
g57034_sb
g57035_da
g57035_db
g57035_sb
g57038_da
g57038_db
g57038_sb
g57039_da
g57039_db
g57039_sb
g57040_da
g57040_db
g57040_sb
g57041_da
g57041_sb
g57042_da
g57042_db
g57042_sb
g57044_da
g57044_db
g57044_sb
g57045_da
g57045_db
g57045_sb
g57046_da
g57046_db
g57046_sb
g57047_da
g57047_db
g57047_sb
g57048_da
g57048_db
g57048_sb
g57049_da
g57049_db
g57049_sb
g57050_da
g57050_db
g57050_sb
g57052_da
g57052_db
g57052_sb
g57053_da
g57053_db
g57053_sb
g57054_da
g57054_db
g57054_sb
g57055_da
g57055_db
g57055_sb
g57056_da
g57056_db
g57056_sb
g57058_da
g57058_db
g57058_sb
g57059_da
g57059_db
g57059_sb
g57060_da
g57060_db
g57060_sb
g57061_da
g57061_db
g57061_sb
g57064_da
g57064_db
g57064_sb
g57065_db
g57068_sb
g57070_da
g57070_db
g57070_sb
g57071_da
g57071_db
g57071_sb
g57072_da
g57072_db
g57072_sb
g57073_da
g57073_db
g57073_sb
g57074_da
g57074_db
g57074_sb
g57075_da
g57075_db
g57075_sb
g57076_da
g57076_db
g57076_sb
g57077_da
g57077_sb
g57078_da
g57078_db
g57078_sb
g57079_da
g57079_db
g57079_sb
g57081_da
g57081_db
g57081_sb
g57082_da
g57082_db
g57082_sb
g57083_da
g57083_db
g57083_sb
g57084_da
g57084_db
g57084_sb
g57085_da
g57085_db
g57085_sb
g57086_da
g57086_db
g57086_sb
g57087_da
g57087_db
g57087_sb
g57088_da
g57088_db
g57088_sb
g57089_da
g57089_db
g57089_sb
g57090_da
g57090_db
g57090_sb
g57091_da
g57091_db
g57091_sb
g57092_da
g57092_db
g57092_sb
g57093_da
g57093_db
g57093_sb
g57095_da
g57095_db
g57095_sb
g57097_da
g57097_db
g57097_sb
g57098_da
g57098_db
g57098_sb
g57099_da
g57099_db
g57099_sb
g57102_da
g57102_db
g57102_sb
g57103_da
g57103_db
g57103_sb
g57105_da
g57105_db
g57105_sb
g57107_da
g57107_db
g57107_sb
g57108_da
g57108_db
g57108_sb
g57109_da
g57109_db
g57109_sb
g57110_da
g57110_db
g57110_sb
g57111_da
g57111_db
g57111_sb
g57112_da
g57112_db
g57112_sb
g57116_da
g57116_db
g57116_sb
g57117_da
g57117_db
g57119_da
g57119_db
g57119_sb
g57120_da
g57120_db
g57120_sb
g57121_da
g57121_db
g57121_sb
g57122_da
g57122_db
g57122_sb
g57123_da
g57123_db
g57123_sb
g57124_da
g57124_db
g57124_sb
g57125_da
g57125_db
g57125_sb
g57126_da
g57126_db
g57126_sb
g57127_da
g57127_db
g57127_sb
g57128_da
g57128_db
g57128_sb
g57130_da
g57130_db
g57130_sb
g57132_da
g57132_db
g57132_sb
g57133_da
g57133_db
g57133_sb
g57134_da
g57134_db
g57134_sb
g57135_da
g57135_db
g57135_sb
g57136_da
g57136_db
g57136_sb
g57137_da
g57137_db
g57137_sb
g57140_da
g57140_db
g57140_sb
g57142_da
g57142_db
g57142_sb
g57143_da
g57143_db
g57143_sb
g57144_da
g57144_db
g57144_sb
g57145_da
g57145_db
g57145_sb
g57147_da
g57147_db
g57147_sb
g57149_sb
g57154_da
g57154_db
g57154_sb
g57155_da
g57155_db
g57156_da
g57156_db
g57156_sb
g57157_da
g57157_db
g57157_sb
g57159_da
g57159_db
g57159_sb
g57160_da
g57160_db
g57160_sb
g57161_da
g57161_db
g57161_sb
g57162_da
g57162_db
g57162_sb
g57163_da
g57163_db
g57163_sb
g57165_da
g57165_db
g57165_sb
g57166_da
g57166_db
g57166_sb
g57167_da
g57167_db
g57168_da
g57168_db
g57168_sb
g57169_da
g57169_db
g57169_sb
g57170_da
g57170_db
g57170_sb
g57171_da
g57171_db
g57171_sb
g57172_da
g57172_db
g57172_sb
g57176_da
g57176_db
g57176_sb
g57179_da
g57179_db
g57179_sb
g57181_da
g57181_db
g57181_sb
g57182_da
g57182_db
g57184_da
g57184_db
g57184_sb
g57185_da
g57185_db
g57185_sb
g57186_da
g57186_db
g57186_sb
g57187_da
g57187_db
g57187_sb
g57188_da
g57188_db
g57188_sb
g57189_da
g57189_db
g57189_sb
g57190_da
g57190_db
g57190_sb
g57192_da
g57192_sb
g57193_da
g57193_db
g57193_sb
g57194_da
g57194_db
g57194_sb
g57195_da
g57195_db
g57195_sb
g57196_db
g57197_da
g57197_db
g57197_sb
g57199_da
g57199_db
g57199_sb
g57200_da
g57200_db
g57200_sb
g57202_da
g57202_db
g57202_sb
g57203_da
g57203_db
g57203_sb
g57205_da
g57205_db
g57205_sb
g57208_da
g57208_db
g57208_sb
g57209_da
g57209_db
g57209_sb
g57210_da
g57210_db
g57210_sb
g57211_da
g57211_db
g57211_sb
g57213_db
g57214_da
g57214_db
g57214_sb
g57215_da
g57215_db
g57215_sb
g57216_da
g57216_db
g57216_sb
g57217_da
g57217_db
g57217_sb
g57218_db
g57219_da
g57219_db
g57219_sb
g57220_da
g57220_db
g57220_sb
g57221_da
g57221_sb
g57222_da
g57222_db
g57222_sb
g57223_da
g57223_db
g57224_da
g57224_db
g57224_sb
g57225_da
g57225_db
g57225_sb
g57227_da
g57227_db
g57227_sb
g57228_da
g57228_db
g57228_sb
g57229_da
g57229_db
g57229_sb
g57230_da
g57230_db
g57230_sb
g57232_da
g57232_db
g57232_sb
g57233_da
g57233_db
g57233_sb
g57234_da
g57234_db
g57234_sb
g57235_da
g57235_db
g57235_sb
g57236_da
g57236_db
g57236_sb
g57237_da
g57237_db
g57239_da
g57239_db
g57239_sb
g57240_da
g57240_db
g57240_sb
g57241_da
g57241_sb
g57242_da
g57242_db
g57242_sb
g57243_da
g57243_db
g57244_da
g57244_db
g57244_sb
g57245_da
g57245_db
g57245_sb
g57247_da
g57247_db
g57247_sb
g57248_da
g57248_db
g57248_sb
g57249_da
g57249_db
g57249_sb
g57250_da
g57250_db
g57250_sb
g57251_da
g57251_db
g57251_sb
g57254_da
g57254_db
g57254_sb
g57255_da
g57255_db
g57255_sb
g57256_da
g57256_db
g57256_sb
g57257_da
g57257_db
g57257_sb
g57258_da
g57258_db
g57258_sb
g57259_da
g57259_db
g57259_sb
g57261_da
g57261_db
g57261_sb
g57262_da
g57262_db
g57262_sb
g57263_da
g57263_db
g57263_sb
g57264_da
g57264_db
g57264_sb
g57265_da
g57265_db
g57265_sb
g57266_da
g57266_db
g57266_sb
g57268_da
g57268_db
g57268_sb
g57269_da
g57269_db
g57271_da
g57271_db
g57271_sb
g57272_da
g57272_db
g57272_sb
g57274_da
g57274_db
g57274_sb
g57275_da
g57275_db
g57275_sb
g57277_da
g57277_db
g57277_sb
g57278_da
g57278_db
g57279_da
g57279_db
g57279_sb
g57280_da
g57280_db
g57280_sb
g57281_da
g57281_db
g57281_sb
g57282_da
g57282_db
g57282_sb
g57283_da
g57283_db
g57283_sb
g57284_da
g57284_db
g57284_sb
g57286_da
g57286_db
g57286_sb
g57288_da
g57288_db
g57288_sb
g57289_da
g57289_db
g57289_sb
g57290_da
g57290_db
g57290_sb
g57291_da
g57291_db
g57291_sb
g57292_da
g57292_db
g57292_sb
g57293_da
g57293_db
g57293_sb
g57294_da
g57294_db
g57294_sb
g57295_da
g57295_db
g57295_sb
g57296_da
g57296_db
g57296_sb
g57298_da
g57298_db
g57298_sb
g57299_da
g57299_db
g57299_sb
g57301_da
g57301_db
g57301_sb
g57303_da
g57303_db
g57303_sb
g57304_da
g57304_db
g57304_sb
g57305_da
g57305_db
g57305_sb
g57306_sb
g57309_da
g57309_db
g57309_sb
g57310_da
g57310_db
g57310_sb
g57311_da
g57311_db
g57311_sb
g57312_da
g57312_db
g57312_sb
g57313_da
g57313_db
g57313_sb
g57314_da
g57314_db
g57314_sb
g57315_da
g57315_db
g57315_sb
g57316_da
g57316_db
g57316_sb
g57317_da
g57317_db
g57317_sb
g57319_da
g57319_db
g57319_sb
g57321_da
g57321_db
g57321_sb
g57322_da
g57322_db
g57322_sb
g57323_da
g57323_db
g57323_sb
g57324_da
g57324_db
g57324_sb
g57325_da
g57325_db
g57325_sb
g57326_da
g57326_db
g57326_sb
g57327_da
g57327_db
g57327_sb
g57328_da
g57328_db
g57328_sb
g57329_da
g57329_db
g57329_sb
g57330_da
g57330_db
g57330_sb
g57331_da
g57331_db
g57331_sb
g57332_da
g57332_db
g57332_sb
g57333_da
g57333_db
g57333_sb
g57335_da
g57335_db
g57335_sb
g57336_da
g57336_db
g57336_sb
g57337_da
g57337_db
g57337_sb
g57338_da
g57338_db
g57338_sb
g57340_da
g57340_db
g57340_sb
g57341_db
g57342_db
g57342_sb
g57343_da
g57343_db
g57343_sb
g57345_da
g57345_db
g57345_sb
g57346_da
g57346_db
g57346_sb
g57347_da
g57347_db
g57347_sb
g57350_da
g57350_db
g57350_sb
g57351_da
g57351_db
g57351_sb
g57352_da
g57352_db
g57352_sb
g57353_da
g57353_sb
g57355_da
g57355_db
g57355_sb
g57356_da
g57356_db
g57356_sb
g57358_da
g57358_db
g57358_sb
g57359_da
g57359_db
g57359_sb
g57360_da
g57360_db
g57360_sb
g57361_da
g57361_db
g57361_sb
g57362_da
g57362_db
g57362_sb
g57364_da
g57364_db
g57364_sb
g57367_da
g57367_db
g57367_sb
g57368_da
g57368_db
g57368_sb
g57370_da
g57370_db
g57371_da
g57371_db
g57371_sb
g57372_da
g57372_db
g57372_sb
g57373_da
g57373_db
g57373_sb
g57374_da
g57374_db
g57374_sb
g57375_da
g57375_db
g57375_sb
g57376_da
g57376_db
g57376_sb
g57377_da
g57377_db
g57377_sb
g57378_da
g57378_db
g57378_sb
g57379_da
g57379_db
g57380_da
g57380_db
g57380_sb
g57381_da
g57381_db
g57381_sb
g57382_da
g57382_db
g57382_sb
g57384_da
g57384_db
g57384_sb
g57386_da
g57386_db
g57386_sb
g57387_da
g57387_db
g57387_sb
g57388_da
g57388_db
g57388_sb
g57389_da
g57389_db
g57389_sb
g57390_da
g57390_db
g57390_sb
g57391_da
g57391_db
g57391_sb
g57392_da
g57392_db
g57392_sb
g57393_da
g57393_db
g57393_sb
g57395_da
g57395_db
g57395_sb
g57396_da
g57396_db
g57396_sb
g57397_da
g57397_db
g57397_sb
g57399_da
g57399_db
g57399_sb
g57401_da
g57401_db
g57401_sb
g57402_da
g57402_db
g57402_sb
g57403_da
g57403_db
g57403_sb
g57404_da
g57404_db
g57404_sb
g57405_da
g57405_db
g57405_sb
g57406_da
g57406_db
g57406_sb
g57407_da
g57407_db
g57409_da
g57409_db
g57409_sb
g57410_da
g57410_db
g57410_sb
g57411_da
g57411_db
g57411_sb
g57412_da
g57412_db
g57412_sb
g57413_da
g57413_db
g57413_sb
g57414_da
g57414_db
g57414_sb
g57415_da
g57415_db
g57415_sb
g57416_da
g57416_db
g57416_sb
g57417_da
g57417_db
g57417_sb
g57418_da
g57418_db
g57418_sb
g57419_da
g57419_db
g57419_sb
g57420_da
g57420_db
g57420_sb
g57421_da
g57421_sb
g57422_da
g57422_db
g57422_sb
g57423_da
g57423_db
g57423_sb
g57424_da
g57424_db
g57424_sb
g57425_da
g57425_db
g57425_sb
g57426_da
g57426_db
g57426_sb
g57427_da
g57427_db
g57427_sb
g57428_da
g57428_db
g57428_sb
g57429_da
g57429_db
g57429_sb
g57432_da
g57432_db
g57432_sb
g57434_da
g57434_db
g57434_sb
g57437_da
g57437_db
g57437_sb
g57439_da
g57439_db
g57439_sb
g57440_da
g57440_db
g57440_sb
g57441_da
g57441_db
g57441_sb
g57442_da
g57442_db
g57442_sb
g57443_da
g57443_db
g57443_sb
g57444_da
g57444_db
g57444_sb
g57447_da
g57447_db
g57447_sb
g57448_da
g57448_db
g57448_sb
g57449_da
g57449_db
g57449_sb
g57450_da
g57450_db
g57450_sb
g57451_da
g57451_db
g57451_sb
g57452_da
g57452_db
g57452_sb
g57453_da
g57453_db
g57453_sb
g57454_da
g57454_db
g57454_sb
g57455_da
g57455_db
g57455_sb
g57456_da
g57456_db
g57456_sb
g57457_da
g57457_db
g57457_sb
g57459_da
g57459_db
g57459_sb
g57460_da
g57460_db
g57460_sb
g57461_da
g57461_db
g57462_da
g57462_db
g57462_sb
g57463_da
g57463_db
g57463_sb
g57464_da
g57464_db
g57464_sb
g57465_da
g57465_db
g57465_sb
g57467_da
g57467_db
g57467_sb
g57468_da
g57468_db
g57468_sb
g57469_da
g57469_db
g57469_sb
g57471_da
g57471_db
g57471_sb
g57473_db
g57475_da
g57475_db
g57475_sb
g57476_da
g57476_db
g57476_sb
g57478_da
g57478_db
g57478_sb
g57481_da
g57481_db
g57481_sb
g57482_da
g57482_db
g57482_sb
g57483_da
g57483_db
g57483_sb
g57484_da
g57484_db
g57484_sb
g57485_da
g57485_db
g57485_sb
g57486_da
g57486_db
g57486_sb
g57487_da
g57487_db
g57487_sb
g57488_da
g57488_db
g57488_sb
g57489_da
g57489_db
g57489_sb
g57490_da
g57490_db
g57490_sb
g57491_da
g57491_db
g57491_sb
g57492_da
g57492_db
g57492_sb
g57493_da
g57493_db
g57493_sb
g57494_da
g57494_db
g57494_sb
g57495_da
g57495_db
g57495_sb
g57497_da
g57497_db
g57497_sb
g57498_da
g57498_db
g57498_sb
g57499_da
g57499_db
g57499_sb
g57500_da
g57500_db
g57500_sb
g57502_da
g57502_db
g57502_sb
g57504_da
g57504_db
g57504_sb
g57506_da
g57506_db
g57506_sb
g57507_da
g57507_db
g57507_sb
g57508_da
g57508_db
g57508_sb
g57510_da
g57510_db
g57510_sb
g57511_da
g57511_db
g57511_sb
g57512_da
g57512_db
g57512_sb
g57513_da
g57513_db
g57513_sb
g57514_da
g57514_db
g57514_sb
g57515_da
g57515_db
g57515_sb
g57516_da
g57516_db
g57516_sb
g57517_da
g57517_db
g57517_sb
g57519_da
g57519_db
g57519_sb
g57520_da
g57520_db
g57520_sb
g57521_da
g57521_db
g57521_sb
g57522_da
g57522_db
g57522_sb
g57523_da
g57523_db
g57523_sb
g57524_da
g57524_db
g57524_sb
g57525_da
g57525_db
g57525_sb
g57526_da
g57526_db
g57526_sb
g57527_da
g57527_db
g57527_sb
g57528_da
g57528_db
g57528_sb
g57529_da
g57529_db
g57529_sb
g57530_da
g57530_db
g57530_sb
g57531_da
g57531_db
g57531_sb
g57532_db
g57532_sb
g57534_da
g57534_db
g57534_sb
g57535_da
g57535_db
g57535_sb
g57536_da
g57536_db
g57536_sb
g57537_da
g57537_db
g57537_sb
g57539_da
g57539_db
g57539_sb
g57540_da
g57540_db
g57540_sb
g57541_da
g57541_db
g57541_sb
g57543_da
g57543_db
g57543_sb
g57544_da
g57544_sb
g57547_da
g57547_db
g57547_sb
g57548_da
g57548_db
g57548_sb
g57553_da
g57553_db
g57553_sb
g57556_da
g57556_db
g57556_sb
g57558_db
g57559_da
g57559_db
g57559_sb
g57561_da
g57561_db
g57561_sb
g57562_da
g57562_db
g57562_sb
g57563_da
g57563_db
g57563_sb
g57568_da
g57568_db
g57568_sb
g57569_da
g57569_db
g57569_sb
g57570_da
g57570_db
g57570_sb
g57571_da
g57571_db
g57571_sb
g57572_da
g57572_db
g57572_sb
g57573_da
g57573_db
g57573_sb
g57574_da
g57574_db
g57574_sb
g57575_da
g57575_db
g57575_sb
g57576_da
g57576_db
g57576_sb
g57577_da
g57577_db
g57577_sb
g57581_da
g57581_db
g57581_sb
g57583_da
g57583_db
g57583_sb
g57584_da
g57584_db
g57584_sb
g57586_da
g57586_db
g57586_sb
g57588_da
g57588_db
g57588_sb
g57589_da
g57589_db
g57589_sb
g57591_da
g57591_db
g57591_sb
g57592_da
g57592_db
g57592_sb
g57595_da
g57595_db
g57595_sb
g57597_da
g57597_db
g57597_sb
g57779_da
g57779_db
g57779_sb
g57780_da
g57780_db
g57780_sb
g57781_da
g57781_db
g57781_sb
g57782_da
g57782_db
g57783_da
g57783_db
g57784_da
g57784_db
g57785_da
g57785_db
g57786_da
g57786_db
g57787_da
g57787_db
g57788_da
g57788_db
g57789_da
g57789_db
g57791_da
g57791_db
g57794_da
g57794_db
g57794_sb
g57795_da
g57795_db
g57796_da
g57796_db
g57797_da
g57797_db
g57798_da
g57798_db
g57798_sb
g57799_da
g57799_db
g57800_da
g57800_db
g57801_da
g57801_db
g57802_da
g57802_db
g57856_p
g57863_p
g57875_da
g57875_db
g57875_sb
g57876_p
g57890_da
g57890_db
g57890_sb
g57891_da
g57891_db
g57891_sb
g57892_da
g57892_db
g57892_sb
g57893_da
g57893_db
g57893_sb
g57895_da
g57895_db
g57895_sb
g57898_da
g57898_db
g57898_sb
g57901_da
g57901_db
g57901_sb
g57902_da
g57902_db
g57902_sb
g57903_da
g57903_db
g57903_sb
g57904_da
g57904_db
g57904_sb
g57906_da
g57906_db
g57906_sb
g57907_da
g57907_db
g57907_sb
g57908_da
g57908_db
g57908_sb
g57909_da
g57909_db
g57910_da
g57910_db
g57910_sb
g57911_da
g57911_db
g57911_sb
g57912_da
g57912_db
g57912_sb
g57913_da
g57913_db
g57913_sb
g57914_da
g57914_db
g57914_sb
g57915_da
g57915_db
g57915_sb
g57918_da
g57918_db
g57918_sb
g57919_da
g57919_db
g57919_sb
g57920_da
g57920_db
g57920_sb
g57921_da
g57921_db
g57921_sb
g57922_da
g57922_db
g57922_sb
g57924_da
g57924_db
g57924_sb
g57925_da
g57925_db
g57925_sb
g57926_da
g57926_db
g57926_sb
g57927_da
g57927_db
g57927_sb
g57928_da
g57928_db
g57928_sb
g57929_da
g57929_db
g57929_sb
g57930_da
g57930_db
g57930_sb
g57932_da
g57932_sb
g57933_da
g57933_db
g57933_sb
g57934_da
g57934_db
g57934_sb
g57935_da
g57935_db
g57935_sb
g57936_da
g57936_db
g57936_sb
g57937_da
g57937_sb
g57938_da
g57938_db
g57938_sb
g57941_da
g57941_db
g57941_sb
g57942_da
g57942_sb
g57944_da
g57944_sb
g57947_da
g57947_db
g57947_sb
g57948_da
g57948_db
g57949_da
g57949_db
g57949_sb
g57950_da
g57950_db
g57950_sb
g57951_da
g57951_db
g57951_sb
g57952_da
g57952_db
g57952_sb
g57953_da
g57953_db
g57953_sb
g57954_da
g57954_db
g57954_sb
g57955_da
g57955_db
g57955_sb
g57956_da
g57956_db
g57956_sb
g57958_da
g57958_db
g57958_sb
g57959_da
g57959_db
g57959_sb
g57960_da
g57960_db
g57960_sb
g57961_da
g57961_db
g57961_sb
g57962_da
g57962_db
g57962_sb
g57963_da
g57963_db
g57963_sb
g57964_da
g57964_db
g57964_sb
g57965_da
g57965_db
g57965_sb
g57966_da
g57966_db
g57966_sb
g57967_da
g57967_db
g57967_sb
g57968_da
g57968_db
g57968_sb
g57969_da
g57969_db
g57969_sb
g57970_da
g57970_db
g57970_sb
g57972_da
g57972_db
g57972_sb
g57973_da
g57973_db
g57973_sb
g57974_da
g57974_db
g57974_sb
g57975_da
g57975_db
g57975_sb
g57976_da
g57976_db
g57976_sb
g57978_da
g57978_db
g57978_sb
g57980_da
g57980_db
g57980_sb
g57981_da
g57981_db
g57981_sb
g57982_da
g57982_db
g57982_sb
g57983_da
g57983_db
g57983_sb
g57984_da
g57984_db
g57984_sb
g57986_da
g57986_db
g57986_sb
g57989_da
g57989_db
g57989_sb
g57992_da
g57992_db
g57992_sb
g57993_da
g57993_db
g57993_sb
g57994_da
g57994_db
g57994_sb
g57995_da
g57995_db
g57995_sb
g57996_da
g57996_db
g57996_sb
g57997_da
g57997_db
g57997_sb
g57999_da
g57999_db
g58000_da
g58000_db
g58000_sb
g58001_da
g58001_db
g58001_sb
g58002_da
g58002_db
g58003_da
g58003_db
g58003_sb
g58004_da
g58004_db
g58004_sb
g58005_da
g58005_db
g58005_sb
g58008_da
g58008_sb
g58009_da
g58009_db
g58009_sb
g58011_da
g58011_db
g58011_sb
g58013_da
g58013_db
g58013_sb
g58014_da
g58014_db
g58014_sb
g58016_da
g58016_db
g58016_sb
g58023_db
g58024_da
g58024_db
g58024_sb
g58025_da
g58025_db
g58025_sb
g58027_da
g58027_db
g58027_sb
g58028_da
g58028_db
g58028_sb
g58030_da
g58030_db
g58030_sb
g58031_da
g58031_db
g58031_sb
g58032_da
g58032_db
g58032_sb
g58033_da
g58033_db
g58033_sb
g58034_da
g58034_db
g58034_sb
g58035_da
g58035_db
g58035_sb
g58036_da
g58036_db
g58036_sb
g58037_da
g58037_db
g58037_sb
g58041_da
g58041_db
g58041_sb
g58044_da
g58044_db
g58044_sb
g58046_da
g58046_db
g58046_sb
g58048_da
g58048_db
g58048_sb
g58049_da
g58049_db
g58050_da
g58050_db
g58050_sb
g58051_da
g58051_db
g58051_sb
g58052_da
g58052_db
g58052_sb
g58053_da
g58053_db
g58053_sb
g58055_da
g58055_db
g58055_sb
g58056_da
g58056_db
g58056_sb
g58057_da
g58057_db
g58057_sb
g58058_sb
g58059_da
g58059_db
g58059_sb
g58060_da
g58060_sb
g58061_da
g58061_db
g58061_sb
g58063_da
g58063_sb
g58064_da
g58064_db
g58066_da
g58066_db
g58067_da
g58067_db
g58067_sb
g58068_da
g58068_db
g58068_sb
g58069_da
g58069_db
g58069_sb
g58070_da
g58070_db
g58070_sb
g58071_da
g58071_db
g58071_sb
g58073_db
g58074_da
g58074_db
g58074_sb
g58075_da
g58075_db
g58075_sb
g58076_da
g58076_db
g58076_sb
g58077_da
g58077_db
g58077_sb
g58079_da
g58079_db
g58079_sb
g58080_da
g58080_db
g58080_sb
g58081_da
g58081_db
g58081_sb
g58082_db
g58083_da
g58083_db
g58083_sb
g58084_da
g58084_db
g58084_sb
g58086_da
g58086_db
g58086_sb
g58087_da
g58087_db
g58087_sb
g58088_da
g58088_db
g58088_sb
g58089_da
g58089_db
g58089_sb
g58091_da
g58091_db
g58091_sb
g58092_da
g58092_db
g58092_sb
g58095_da
g58095_db
g58095_sb
g58096_da
g58096_db
g58096_sb
g58099_da
g58099_db
g58099_sb
g58100_da
g58100_db
g58100_sb
g58102_da
g58102_db
g58102_sb
g58103_da
g58103_db
g58103_sb
g58106_da
g58106_db
g58106_sb
g58107_da
g58107_db
g58109_da
g58109_db
g58110_da
g58110_db
g58110_sb
g58111_da
g58111_db
g58111_sb
g58112_da
g58112_db
g58112_sb
g58113_da
g58113_db
g58113_sb
g58116_da
g58116_db
g58116_sb
g58117_da
g58117_db
g58117_sb
g58118_da
g58118_db
g58118_sb
g58119_da
g58119_db
g58119_sb
g58120_da
g58120_db
g58120_sb
g58121_da
g58121_db
g58121_sb
g58123_da
g58123_db
g58124_da
g58124_db
g58124_sb
g58125_da
g58125_db
g58125_sb
g58126_da
g58126_db
g58126_sb
g58127_da
g58127_db
g58127_sb
g58128_da
g58128_db
g58128_sb
g58129_da
g58129_db
g58129_sb
g58130_da
g58130_db
g58130_sb
g58133_da
g58133_db
g58133_sb
g58134_da
g58134_db
g58136_da
g58136_db
g58136_sb
g58137_da
g58137_db
g58137_sb
g58139_da
g58139_db
g58139_sb
g58140_db
g58141_da
g58141_db
g58141_sb
g58142_da
g58142_db
g58142_sb
g58143_da
g58143_db
g58143_sb
g58144_da
g58144_db
g58144_sb
g58145_da
g58145_db
g58145_sb
g58146_da
g58146_db
g58146_sb
g58148_da
g58148_db
g58148_sb
g58150_da
g58150_db
g58150_sb
g58151_da
g58151_db
g58151_sb
g58152_da
g58152_db
g58152_sb
g58153_da
g58153_db
g58153_sb
g58154_db
g58155_da
g58155_db
g58155_sb
g58156_da
g58156_db
g58156_sb
g58157_da
g58157_db
g58157_sb
g58158_da
g58158_db
g58158_sb
g58160_da
g58160_db
g58162_da
g58162_db
g58162_sb
g58163_da
g58163_db
g58163_sb
g58165_da
g58165_db
g58165_sb
g58166_da
g58166_db
g58166_sb
g58167_da
g58167_db
g58167_sb
g58170_da
g58170_db
g58170_sb
g58171_db
g58172_da
g58172_db
g58172_sb
g58173_da
g58173_db
g58173_sb
g58174_da
g58174_db
g58174_sb
g58175_da
g58175_db
g58175_sb
g58176_da
g58176_db
g58176_sb
g58178_da
g58178_db
g58178_sb
g58180_da
g58180_db
g58180_sb
g58181_da
g58181_db
g58181_sb
g58182_da
g58182_db
g58182_sb
g58183_da
g58183_db
g58183_sb
g58184_da
g58184_db
g58184_sb
g58185_da
g58185_db
g58185_sb
g58186_da
g58186_db
g58186_sb
g58187_da
g58187_db
g58187_sb
g58188_da
g58188_db
g58188_sb
g58189_da
g58189_db
g58191_da
g58191_db
g58191_sb
g58192_da
g58192_db
g58192_sb
g58193_da
g58193_db
g58193_sb
g58194_da
g58194_db
g58194_sb
g58195_da
g58195_db
g58195_sb
g58196_da
g58196_db
g58196_sb
g58198_da
g58198_db
g58198_sb
g58199_da
g58199_db
g58200_da
g58200_db
g58200_sb
g58202_da
g58202_db
g58202_sb
g58203_da
g58203_db
g58203_sb
g58204_da
g58204_db
g58204_sb
g58207_da
g58207_db
g58207_sb
g58208_da
g58208_db
g58208_sb
g58209_da
g58209_db
g58209_sb
g58210_da
g58210_db
g58210_sb
g58212_da
g58212_db
g58212_sb
g58213_da
g58213_db
g58215_da
g58215_db
g58215_sb
g58216_da
g58216_db
g58216_sb
g58217_da
g58217_db
g58217_sb
g58218_da
g58218_db
g58218_sb
g58219_da
g58219_db
g58219_sb
g58221_da
g58221_db
g58221_sb
g58224_da
g58224_db
g58224_sb
g58225_da
g58225_db
g58225_sb
g58228_da
g58228_db
g58228_sb
g58229_da
g58229_db
g58229_sb
g58230_da
g58230_db
g58230_sb
g58231_da
g58231_db
g58231_sb
g58232_da
g58232_db
g58232_sb
g58233_da
g58233_db
g58233_sb
g58234_da
g58234_db
g58234_sb
g58235_da
g58235_db
g58235_sb
g58236_da
g58236_db
g58236_sb
g58237_da
g58237_db
g58237_sb
g58238_da
g58238_db
g58238_sb
g58239_da
g58239_db
g58239_sb
g58240_da
g58240_db
g58240_sb
g58241_da
g58241_db
g58241_sb
g58243_da
g58243_db
g58243_sb
g58244_da
g58244_db
g58244_sb
g58245_da
g58245_db
g58245_sb
g58246_da
g58246_db
g58246_sb
g58247_da
g58247_db
g58247_sb
g58248_da
g58248_db
g58248_sb
g58249_da
g58249_db
g58249_sb
g58250_da
g58250_db
g58250_sb
g58252_da
g58252_db
g58252_sb
g58253_da
g58253_db
g58253_sb
g58255_da
g58255_db
g58255_sb
g58257_da
g58257_db
g58257_sb
g58258_da
g58258_db
g58258_sb
g58259_da
g58259_db
g58259_sb
g58260_da
g58260_db
g58260_sb
g58261_da
g58261_db
g58261_sb
g58265_da
g58265_db
g58266_da
g58266_db
g58266_sb
g58268_da
g58268_db
g58268_sb
g58269_da
g58269_db
g58269_sb
g58272_da
g58272_db
g58272_sb
g58273_da
g58273_db
g58273_sb
g58274_da
g58274_db
g58274_sb
g58275_da
g58275_db
g58275_sb
g58276_da
g58276_db
g58276_sb
g58277_da
g58277_db
g58277_sb
g58278_da
g58278_db
g58278_sb
g58279_da
g58279_db
g58279_sb
g58280_da
g58280_db
g58280_sb
g58281_da
g58281_db
g58281_sb
g58282_da
g58282_db
g58282_sb
g58283_da
g58283_db
g58283_sb
g58285_da
g58285_db
g58285_sb
g58286_da
g58286_db
g58286_sb
g58287_da
g58287_db
g58287_sb
g58288_da
g58288_db
g58288_sb
g58289_da
g58289_db
g58289_sb
g58290_da
g58290_db
g58290_sb
g58291_da
g58291_db
g58291_sb
g58292_da
g58292_db
g58292_sb
g58295_da
g58295_db
g58295_sb
g58297_da
g58297_db
g58297_sb
g58299_db
g58300_da
g58300_db
g58300_sb
g58302_da
g58302_db
g58302_sb
g58303_da
g58303_db
g58303_sb
g58304_da
g58304_db
g58304_sb
g58305_da
g58305_db
g58305_sb
g58306_da
g58306_db
g58306_sb
g58307_da
g58307_db
g58307_sb
g58310_da
g58310_db
g58310_sb
g58311_da
g58311_db
g58311_sb
g58312_da
g58312_db
g58312_sb
g58313_da
g58313_db
g58313_sb
g58314_da
g58314_sb
g58315_da
g58315_db
g58315_sb
g58316_da
g58316_db
g58316_sb
g58317_da
g58317_db
g58317_sb
g58318_da
g58318_db
g58318_sb
g58319_da
g58319_db
g58319_sb
g58321_da
g58321_db
g58321_sb
g58322_da
g58322_sb
g58323_da
g58323_db
g58323_sb
g58324_da
g58324_db
g58324_sb
g58325_da
g58325_db
g58325_sb
g58326_da
g58326_db
g58326_sb
g58327_da
g58327_db
g58327_sb
g58328_da
g58328_db
g58328_sb
g58329_da
g58329_db
g58329_sb
g58330_da
g58330_db
g58330_sb
g58332_da
g58332_db
g58332_sb
g58333_da
g58333_db
g58333_sb
g58336_da
g58336_db
g58336_sb
g58337_da
g58337_db
g58337_sb
g58339_da
g58339_db
g58341_sb
g58342_da
g58342_db
g58342_sb
g58343_da
g58343_db
g58343_sb
g58344_da
g58344_db
g58344_sb
g58345_da
g58345_db
g58345_sb
g58346_da
g58346_db
g58346_sb
g58347_da
g58347_db
g58347_sb
g58348_da
g58348_db
g58348_sb
g58349_da
g58349_db
g58349_sb
g58350_da
g58350_db
g58350_sb
g58351_da
g58351_db
g58351_sb
g58352_da
g58352_db
g58352_sb
g58353_da
g58353_db
g58353_sb
g58354_da
g58354_db
g58354_sb
g58355_da
g58355_sb
g58357_da
g58357_db
g58357_sb
g58358_da
g58358_db
g58358_sb
g58359_da
g58359_db
g58359_sb
g58360_da
g58360_db
g58360_sb
g58361_da
g58361_sb
g58362_da
g58362_db
g58362_sb
g58363_da
g58363_db
g58363_sb
g58364_da
g58364_db
g58364_sb
g58366_da
g58366_db
g58366_sb
g58367_da
g58367_db
g58367_sb
g58369_da
g58369_db
g58369_sb
g58370_da
g58370_db
g58370_sb
g58371_da
g58371_db
g58371_sb
g58372_da
g58372_db
g58372_sb
g58373_da
g58373_db
g58373_sb
g58374_da
g58374_db
g58374_sb
g58375_da
g58375_db
g58375_sb
g58376_da
g58376_db
g58376_sb
g58378_da
g58378_db
g58378_sb
g58379_da
g58379_db
g58379_sb
g58380_da
g58380_db
g58380_sb
g58381_da
g58381_db
g58381_sb
g58382_da
g58382_db
g58382_sb
g58383_da
g58383_sb
g58384_da
g58384_db
g58384_sb
g58385_da
g58385_db
g58385_sb
g58386_da
g58386_db
g58386_sb
g58387_da
g58387_db
g58387_sb
g58388_da
g58388_db
g58388_sb
g58389_da
g58389_db
g58389_sb
g58390_da
g58390_db
g58390_sb
g58393_da
g58393_sb
g58394_da
g58394_db
g58394_sb
g58395_da
g58395_db
g58395_sb
g58397_da
g58397_db
g58397_sb
g58398_da
g58398_db
g58398_sb
g58399_da
g58399_db
g58399_sb
g58401_da
g58401_db
g58401_sb
g58402_db
g58404_da
g58404_db
g58404_sb
g58405_da
g58405_db
g58405_sb
g58406_da
g58406_db
g58406_sb
g58409_da
g58409_db
g58409_sb
g58411_da
g58411_db
g58411_sb
g58413_da
g58413_db
g58413_sb
g58415_da
g58415_db
g58415_sb
g58416_da
g58416_db
g58416_sb
g58419_da
g58419_db
g58419_sb
g58421_da
g58421_db
g58421_sb
g58425_da
g58425_db
g58425_sb
g58426_da
g58426_db
g58427_da
g58427_db
g58427_sb
g58428_da
g58428_sb
g58429_da
g58429_db
g58429_sb
g58430_da
g58430_db
g58430_sb
g58431_da
g58431_db
g58431_sb
g58433_db
g58434_da
g58434_db
g58436_da
g58436_db
g58436_sb
g58437_da
g58437_db
g58438_db
g58439_da
g58439_db
g58439_sb
g58440_da
g58440_db
g58440_sb
g58441_da
g58441_db
g58441_sb
g58442_da
g58442_db
g58442_sb
g58443_da
g58443_db
g58443_sb
g58445_da
g58445_db
g58445_sb
g58447_da
g58447_db
g58447_sb
g58448_da
g58448_db
g58448_sb
g58449_da
g58449_db
g58449_sb
g58450_da
g58450_db
g58450_sb
g58453_da
g58453_db
g58453_sb
g58455_da
g58455_db
g58455_sb
g58456_da
g58456_db
g58456_sb
g58457_da
g58457_db
g58457_sb
g58459_da
g58459_db
g58459_sb
g58460_da
g58460_db
g58460_sb
g58461_da
g58461_db
g58461_sb
g58462_da
g58462_db
g58462_sb
g58463_da
g58463_db
g58463_sb
g58464_da
g58464_db
g58464_sb
g58465_da
g58465_db
g58465_sb
g58466_da
g58466_db
g58466_sb
g58467_da
g58467_db
g58467_sb
g58468_da
g58468_db
g58468_sb
g58469_da
g58469_db
g58469_sb
g58470_da
g58470_db
g58470_sb
g58471_da
g58471_db
g58471_sb
g58472_da
g58472_db
g58472_sb
g58473_da
g58473_db
g58473_sb
g58474_da
g58474_db
g58474_sb
g58475_da
g58475_db
g58475_sb
g58476_da
g58476_db
g58476_sb
g58477_da
g58477_db
g58477_sb
g58478_da
g58478_db
g58478_sb
g58479_da
g58479_db
g58479_sb
g58480_da
g58480_db
g58480_sb
g58481_da
g58481_db
g58481_sb
g58483_da
g58483_db
g58483_sb
g58484_da
g58484_db
g58484_sb
g58485_da
g58485_db
g58485_sb
g58486_da
g58486_db
g58486_sb
g58487_da
g58487_db
g58487_sb
g58488_da
g58488_db
g58488_sb
g58489_da
g58489_db
g58489_sb
g58490_p
g58569_p
g58576_da
g58576_db
g58582_p
g58590_da
g58590_db
g58590_sb
g58591_da
g58591_db
g58597_da
g58597_db
g58597_sb
g58598_da
g58598_db
g58598_sb
g58599_p
g58600_da
g58600_db
g58600_sb
g58601_da
g58601_db
g58601_sb
g58605_da
g58605_db
g58605_sb
g58606_da
g58606_db
g58608_da
g58608_db
g58608_sb
g58610_da
g58610_db
g58610_sb
g58616_da
g58616_db
g58616_sb
g58617_da
g58617_db
g58617_sb
g58618_da
g58618_db
g58618_sb
g58619_da
g58619_db
g58619_sb
g58620_da
g58620_db
g58620_sb
g58621_da
g58621_db
g58621_sb
g58622_da
g58622_db
g58622_sb
g58630_da
g58630_db
g58630_sb
g58631_da
g58631_db
g58631_sb
g58632_da
g58632_db
g58632_sb
g58633_da
g58633_db
g58633_sb
g58634_da
g58634_db
g58634_sb
g58635_da
g58635_db
g58635_sb
g58636_da
g58636_db
g58636_sb
g58640_da
g58640_db
g58640_sb
g58652_da
g58652_db
g58652_sb
g58653_da
g58653_db
g58653_sb
g58654_da
g58654_db
g58654_sb
g58655_da
g58655_db
g58655_sb
g58692_p
g58695_p
g58742_p
g58744_p
g58759_p
g58760_p
g58761_p
g58763_p
g58764_p
g58767_da
g58767_db
g58767_sb
g58768_da
g58768_db
g58768_sb
g58769_da
g58769_db
g58769_sb
g58770_da
g58770_db
g58770_sb
g58771_da
g58771_db
g58771_sb
g58772_da
g58772_db
g58772_sb
g58773_da
g58773_db
g58773_sb
g58774_da
g58774_db
g58774_sb
g58775_da
g58775_db
g58775_sb
g58776_da
g58776_db
g58776_sb
g58777_da
g58777_db
g58777_sb
g58778_da
g58778_db
g58778_sb
g58779_da
g58779_db
g58779_sb
g58780_da
g58780_db
g58780_sb
g58781_da
g58781_db
g58781_sb
g58782_da
g58782_db
g58782_sb
g58783_da
g58783_db
g58783_sb
g58784_da
g58784_db
g58784_sb
g58785_da
g58785_db
g58785_sb
g58786_da
g58786_db
g58786_sb
g58787_da
g58787_db
g58787_sb
g58788_da
g58788_db
g58788_sb
g58789_da
g58789_db
g58789_sb
g58790_da
g58790_db
g58790_sb
g58791_da
g58791_db
g58791_sb
g58792_da
g58792_db
g58792_sb
g58793_da
g58793_db
g58793_sb
g58795_da
g58795_db
g58795_sb
g58796_da
g58796_db
g58796_sb
g58797_da
g58797_db
g58797_sb
g58798_da
g58798_db
g58798_sb
g58799_da
g58799_db
g58799_sb
g58800_da
g58800_db
g58800_sb
g58801_da
g58801_db
g58801_sb
g58802_da
g58802_db
g58802_sb
g58803_da
g58803_db
g58803_sb
g58804_da
g58804_db
g58804_sb
g58805_da
g58805_db
g58805_sb
g58806_da
g58806_db
g58806_sb
g58807_da
g58807_db
g58807_sb
g58808_da
g58808_db
g58808_sb
g58809_da
g58809_db
g58809_sb
g58810_da
g58810_db
g58810_sb
g58811_da
g58811_db
g58811_sb
g58812_da
g58812_db
g58812_sb
g58813_da
g58813_db
g58813_sb
g58814_da
g58814_db
g58814_sb
g58815_da
g58815_db
g58815_sb
g58816_da
g58816_db
g58816_sb
g58817_da
g58817_db
g58817_sb
g58818_da
g58818_db
g58818_sb
g58819_da
g58819_db
g58819_sb
g58820_da
g58820_db
g58820_sb
g58821_da
g58821_db
g58821_sb
g58822_da
g58822_db
g58822_sb
g58823_da
g58823_db
g58823_sb
g58824_da
g58824_db
g58824_sb
g58825_da
g58825_db
g58825_sb
g58829_db
g58830_da
g58830_db
g58830_sb
g58831_da
g58831_db
g58831_sb
g58832_da
g58832_db
g58833_da
g58833_db
g58833_sb
g58834_da
g58834_db
g58834_sb
g58835_da
g58835_db
g58835_sb
g58836_da
g58836_db
g58836_sb
g58840_da
g58840_db
g58840_sb
g58842_da
g58842_db
g58842_sb
g58843_da
g58843_db
g58843_sb
g59082_da
g59082_db
g59082_sb
g59086_p
g59089_da
g59089_db
g59089_sb
g59090_da
g59090_db
g59090_sb
g59091_da
g59091_db
g59091_sb
g59095_p
g59096_da
g59096_db
g59096_sb
g59098_da
g59098_db
g59098_sb
g59109_da
g59109_db
g59109_sb
g59110_da
g59110_db
g59110_sb
g59111_da
g59111_db
g59111_sb
g59112_da
g59112_db
g59112_sb
g59113_da
g59113_db
g59113_sb
g59114_da
g59114_db
g59114_sb
g59115_da
g59115_db
g59115_sb
g59116_da
g59116_db
g59116_sb
g59117_da
g59117_db
g59117_sb
g59118_da
g59118_db
g59118_sb
g59119_da
g59119_db
g59119_sb
g59120_da
g59120_db
g59120_sb
g59121_da
g59121_db
g59121_sb
g59122_da
g59122_db
g59122_sb
g59123_da
g59123_db
g59123_sb
g59124_p
g59125_p
g59127_p
g59128_p
g59196_p
g59198_p
g59199_p
g59201_p
g59227_p
g59228_p
g59229_p
g59230_da
g59230_db
g59230_sb
g59231_da
g59231_db
g59231_sb
g59232_AP
g59232_BP
g59232_p
g59234_da
g59234_db
g59234_sb
g59240_da
g59240_db
g59240_sb
g59300_p
g59331_p
g59343_p
g59344_p
g59346_p
g59347_p
g59350_da
g59350_db
g59350_sb
g59364_p
g59368_da
g59368_db
g59368_sb
g59369_da
g59369_db
g59369_sb
g59370_da
g59370_db
g59370_sb
g59371_da
g59371_db
g59371_sb
g59372_da
g59372_db
g59372_sb
g59373_da
g59373_db
g59373_sb
g59374_p
g59378_da
g59378_db
g59378_sb
g59379_da
g59379_db
g59379_sb
g59380_da
g59380_db
g59380_sb
g59381_da
g59381_db
g59381_sb
g59382_da
g59382_db
g59382_sb
g59383_da
g59383_db
g59383_sb
g59384_sb
g59385_p
g59386_p
g59387_da
g59387_db
g59387_sb
g59388_p
g59389_p
g59622_p
g59623_p
g59627_p
g59659_p
g59665_p
g59666_p
g59670_p
g59674_p
g59721_p
g59761_p
g59770_da
g59770_db
g59783_p
g59790_p
g59791_p
g59793_p
g59794_p
g59795_p
g59797_da
g59797_db
g59797_sb
g59798_da
g59798_db
g59798_sb
g59800_da
g59800_db
g59800_sb
g59801_da
g59801_db
g59801_sb
g59802_p
g59803_p
g59804_da
g59804_db
g59804_sb
g59805_da
g59805_db
g59805_sb
g59806_da
g59806_db
g59806_sb
g59807_da
g59807_db
g59807_sb
g59808_da
g59808_db
g59808_sb
g59809_da
g59809_db
g59809_sb
g60298_p
g60304_p
g60307_p
g60310_p
g60319_p
g60330_p
g60408_db
g60414_p
g60415_p
g60557_p
g60591_p
g60604_da
g60604_sb
g60605_da
g60605_sb
g60606_da
g60606_db
g60606_sb
g60607_da
g60607_db
g60607_sb
g60608_da
g60608_db
g60608_sb
g60609_da
g60609_db
g60609_sb
g60610_da
g60610_db
g60610_sb
g60611_da
g60611_db
g60611_sb
g60612_da
g60612_db
g60612_sb
g60613_da
g60613_db
g60613_sb
g60614_da
g60614_sb
g60615_db
g60616_da
g60616_db
g60616_sb
g60617_da
g60617_db
g60617_sb
g60618_da
g60618_db
g60618_sb
g60619_da
g60619_sb
g60620_da
g60620_db
g60620_sb
g60621_da
g60621_db
g60621_sb
g60622_da
g60622_db
g60622_sb
g60623_da
g60623_db
g60623_sb
g60624_da
g60624_db
g60624_sb
g60625_da
g60625_db
g60625_sb
g60626_da
g60626_db
g60626_sb
g60627_da
g60627_db
g60627_sb
g60628_da
g60628_db
g60628_sb
g60629_da
g60629_db
g60629_sb
g60630_da
g60630_sb
g60631_da
g60631_db
g60631_sb
g60633_da
g60633_db
g60633_sb
g60634_da
g60634_db
g60634_sb
g60635_da
g60635_sb
g60636_da
g60636_db
g60636_sb
g60637_da
g60637_db
g60637_sb
g60638_da
g60638_db
g60638_sb
g60639_da
g60639_db
g60639_sb
g60640_da
g60640_db
g60640_sb
g60641_da
g60641_db
g60641_sb
g60642_da
g60642_sb
g60643_da
g60643_db
g60643_sb
g60644_da
g60644_db
g60644_sb
g60645_da
g60645_db
g60645_sb
g60646_da
g60646_db
g60646_sb
g60647_da
g60647_db
g60647_sb
g60648_da
g60648_db
g60648_sb
g60649_da
g60649_db
g60649_sb
g60650_da
g60650_db
g60650_sb
g60651_da
g60651_db
g60651_sb
g60652_da
g60652_db
g60652_sb
g60653_da
g60653_db
g60653_sb
g60654_da
g60654_sb
g60655_da
g60655_db
g60655_sb
g60656_da
g60656_db
g60656_sb
g60657_da
g60657_sb
g60658_da
g60658_db
g60658_sb
g60659_sb
g60660_da
g60660_db
g60660_sb
g60661_da
g60661_db
g60661_sb
g60662_da
g60662_db
g60662_sb
g60664_da
g60664_db
g60664_sb
g60666_da
g60666_db
g60667_da
g60667_db
g60667_sb
g60668_da
g60668_sb
g60669_da
g60669_db
g60669_sb
g60670_da
g60670_db
g60670_sb
g60673_da
g60673_sb
g60675_da
g60675_db
g60675_sb
g60676_da
g60676_db
g60676_sb
g60677_da
g60677_db
g60677_sb
g60678_da
g60678_db
g60678_sb
g60679_da
g60679_db
g60679_sb
g60681_da
g60681_db
g60681_sb
g60682_da
g60682_db
g60686_da
g60686_db
g60686_sb
g60687_da
g60687_db
g60687_sb
g60688_da
g60688_db
g60688_sb
g60689_da
g60689_db
g60689_sb
g60691_da
g60691_db
g60691_sb
g60692_da
g60692_db
g60692_sb
g60693_p
g60694_p
g60695_p
g60696_p
g60698_p
g61569_p
g61570_p
g61575_p
g61597_p
g61606_p
g61618_AP
g61618_BP
g61618_p
g61622_p
g61636_p
g61637_p
g61654_p
g61676_da
g61676_db
g61676_sb
g61689_p
g61693_p
g61697_da
g61697_db
g61697_sb
g61699_da
g61699_db
g61699_sb
g61701_da
g61701_db
g61701_sb
g61702_da
g61702_db
g61702_sb
g61703_da
g61703_db
g61703_sb
g61704_da
g61704_db
g61704_sb
g61705_da
g61705_db
g61705_sb
g61706_da
g61706_db
g61706_sb
g61707_da
g61707_db
g61707_sb
g61708_da
g61708_db
g61708_sb
g61709_da
g61709_db
g61709_sb
g61710_da
g61710_db
g61710_sb
g61711_da
g61711_db
g61711_sb
g61712_da
g61712_db
g61712_sb
g61713_da
g61713_db
g61713_sb
g61714_da
g61714_db
g61714_sb
g61715_da
g61715_db
g61715_sb
g61716_da
g61716_db
g61716_sb
g61717_da
g61717_db
g61717_sb
g61720_da
g61720_db
g61720_sb
g61721_da
g61721_db
g61721_sb
g61724_da
g61724_db
g61724_sb
g61725_da
g61725_db
g61725_sb
g61726_da
g61726_db
g61726_sb
g61727_da
g61727_db
g61727_sb
g61728_da
g61728_db
g61728_sb
g61730_da
g61730_db
g61730_sb
g61731_da
g61731_db
g61731_sb
g61732_da
g61732_db
g61732_sb
g61733_da
g61733_db
g61734_da
g61734_db
g61734_sb
g61735_da
g61735_db
g61735_sb
g61736_da
g61736_db
g61736_sb
g61737_da
g61737_db
g61737_sb
g61738_da
g61738_db
g61738_sb
g61739_da
g61739_db
g61739_sb
g61740_da
g61740_db
g61740_sb
g61741_da
g61741_db
g61741_sb
g61742_da
g61742_db
g61742_sb
g61743_da
g61743_db
g61743_sb
g61744_da
g61744_db
g61744_sb
g61745_da
g61745_db
g61745_sb
g61746_da
g61746_db
g61746_sb
g61747_da
g61747_db
g61747_sb
g61748_da
g61748_db
g61748_sb
g61749_da
g61749_db
g61749_sb
g61750_da
g61750_db
g61750_sb
g61753_da
g61753_db
g61753_sb
g61754_da
g61754_db
g61754_sb
g61755_da
g61755_db
g61755_sb
g61757_da
g61757_db
g61757_sb
g61759_da
g61759_db
g61759_sb
g61760_da
g61760_db
g61760_sb
g61761_da
g61761_db
g61761_sb
g61763_da
g61763_db
g61763_sb
g61764_da
g61764_db
g61764_sb
g61765_da
g61765_db
g61765_sb
g61767_da
g61767_db
g61767_sb
g61768_da
g61768_db
g61768_sb
g61769_da
g61769_db
g61769_sb
g61770_da
g61770_db
g61770_sb
g61771_da
g61771_db
g61771_sb
g61772_da
g61772_db
g61772_sb
g61773_da
g61773_db
g61773_sb
g61774_da
g61774_db
g61774_sb
g61775_da
g61775_db
g61775_sb
g61776_da
g61776_db
g61776_sb
g61777_da
g61777_db
g61777_sb
g61778_da
g61778_db
g61778_sb
g61779_da
g61779_db
g61779_sb
g61781_da
g61781_db
g61781_sb
g61782_da
g61782_db
g61782_sb
g61783_da
g61783_db
g61783_sb
g61787_da
g61787_db
g61787_sb
g61790_da
g61790_db
g61790_sb
g61792_da
g61792_db
g61792_sb
g61793_da
g61793_db
g61794_da
g61794_db
g61794_sb
g61796_da
g61796_db
g61796_sb
g61797_da
g61797_db
g61797_sb
g61798_da
g61798_db
g61798_sb
g61800_da
g61800_db
g61800_sb
g61801_da
g61801_db
g61801_sb
g61802_da
g61802_db
g61802_sb
g61803_da
g61803_db
g61803_sb
g61804_da
g61804_db
g61804_sb
g61805_da
g61805_db
g61805_sb
g61806_da
g61806_db
g61806_sb
g61807_da
g61807_db
g61807_sb
g61808_da
g61808_db
g61808_sb
g61809_da
g61809_db
g61809_sb
g61810_da
g61810_db
g61810_sb
g61811_da
g61811_db
g61811_sb
g61812_da
g61812_db
g61812_sb
g61814_da
g61814_db
g61814_sb
g61815_da
g61815_db
g61815_sb
g61816_da
g61816_db
g61816_sb
g61820_da
g61820_db
g61820_sb
g61823_da
g61823_db
g61823_sb
g61824_da
g61824_db
g61824_sb
g61825_da
g61825_db
g61825_sb
g61826_da
g61826_db
g61826_sb
g61827_da
g61827_db
g61827_sb
g61829_da
g61829_db
g61829_sb
g61830_da
g61830_sb
g61832_p
g61833_p
g61834_p
g61838_p
g61839_p
g61840_da
g61840_db
g61840_sb
g61846_p
g61850_p
g61851_p
g61855_da
g61855_db
g61855_sb
g61856_da
g61856_db
g61856_sb
g61857_p
g61858_da
g61858_db
g61858_sb
g61859_da
g61859_db
g61859_sb
g61860_da
g61860_db
g61861_da
g61861_db
g61861_sb
g61862_da
g61862_db
g61862_sb
g61863_da
g61863_db
g61863_sb
g61864_da
g61864_db
g61864_sb
g61865_da
g61865_db
g61865_sb
g61866_da
g61866_sb
g61868_da
g61868_db
g61868_sb
g61869_da
g61869_db
g61869_sb
g61870_da
g61870_db
g61870_sb
g61873_da
g61873_db
g61873_sb
g61874_da
g61874_db
g61874_sb
g61875_da
g61875_db
g61877_da
g61877_db
g61877_sb
g61878_da
g61878_db
g61878_sb
g61879_da
g61879_db
g61879_sb
g61880_da
g61880_db
g61880_sb
g61881_da
g61881_db
g61881_sb
g61885_da
g61885_db
g61885_sb
g61886_da
g61886_db
g61886_sb
g61887_da
g61887_db
g61887_sb
g61889_da
g61889_db
g61889_sb
g61890_da
g61890_db
g61890_sb
g61891_da
g61891_db
g61891_sb
g61892_da
g61892_db
g61892_sb
g61893_da
g61893_db
g61893_sb
g61894_da
g61894_db
g61894_sb
g61895_da
g61895_db
g61895_sb
g61896_da
g61896_db
g61896_sb
g61897_da
g61897_db
g61897_sb
g61898_da
g61898_db
g61898_sb
g61899_da
g61899_db
g61899_sb
g61900_da
g61900_db
g61900_sb
g61901_da
g61901_db
g61901_sb
g61903_da
g61903_db
g61903_sb
g61904_da
g61904_db
g61904_sb
g61905_da
g61905_db
g61905_sb
g61908_da
g61908_db
g61908_sb
g61910_da
g61910_db
g61910_sb
g61912_da
g61912_db
g61912_sb
g61913_da
g61913_db
g61913_sb
g61914_da
g61914_db
g61914_sb
g61915_da
g61915_db
g61915_sb
g61916_da
g61916_db
g61916_sb
g61918_da
g61918_db
g61918_sb
g61920_da
g61920_db
g61920_sb
g61922_da
g61922_db
g61922_sb
g61923_da
g61923_db
g61923_sb
g61924_da
g61924_db
g61924_sb
g61925_da
g61925_db
g61925_sb
g61926_da
g61926_db
g61926_sb
g61927_da
g61927_db
g61927_sb
g61928_da
g61928_db
g61928_sb
g61929_da
g61929_db
g61929_sb
g61930_da
g61930_db
g61930_sb
g61931_da
g61931_db
g61931_sb
g61932_da
g61932_db
g61932_sb
g61933_da
g61933_db
g61933_sb
g61934_da
g61934_db
g61934_sb
g61935_da
g61935_db
g61935_sb
g61937_da
g61937_db
g61937_sb
g61938_da
g61938_db
g61938_sb
g61939_da
g61939_db
g61939_sb
g61942_da
g61942_db
g61942_sb
g61943_da
g61943_db
g61943_sb
g61945_da
g61945_db
g61945_sb
g61946_da
g61946_sb
g61947_da
g61947_db
g61947_sb
g61949_da
g61949_db
g61949_sb
g61950_da
g61950_db
g61950_sb
g61951_da
g61951_db
g61951_sb
g61953_da
g61953_db
g61953_sb
g61954_da
g61954_db
g61954_sb
g61958_da
g61958_db
g61958_sb
g61959_da
g61959_db
g61959_sb
g61960_da
g61960_db
g61960_sb
g61961_da
g61961_db
g61961_sb
g61962_da
g61962_db
g61962_sb
g61964_da
g61964_db
g61964_sb
g61965_da
g61965_db
g61966_da
g61966_db
g61966_sb
g61967_da
g61967_db
g61967_sb
g61968_da
g61968_db
g61968_sb
g61969_da
g61969_db
g61969_sb
g61970_da
g61970_db
g61970_sb
g61971_da
g61971_db
g61971_sb
g61972_da
g61972_db
g61972_sb
g61973_da
g61973_db
g61973_sb
g61974_da
g61974_db
g61974_sb
g61975_da
g61975_db
g61975_sb
g61976_da
g61976_db
g61976_sb
g61977_da
g61977_db
g61977_sb
g61978_da
g61978_db
g61978_sb
g61979_da
g61979_db
g61979_sb
g61980_da
g61980_db
g61980_sb
g61981_da
g61981_db
g61981_sb
g61982_da
g61982_db
g61982_sb
g61983_da
g61983_db
g61983_sb
g61984_da
g61984_db
g61984_sb
g61985_da
g61985_db
g61985_sb
g61986_da
g61986_db
g61986_sb
g61987_da
g61987_db
g61987_sb
g61988_da
g61988_db
g61988_sb
g61989_da
g61989_db
g61989_sb
g61990_da
g61990_db
g61990_sb
g61992_da
g61992_db
g61992_sb
g61993_da
g61993_db
g61993_sb
g61994_da
g61994_db
g61994_sb
g61995_da
g61995_db
g61995_sb
g61996_da
g61996_db
g61996_sb
g61997_da
g61997_db
g61997_sb
g61998_da
g61998_db
g61998_sb
g61999_da
g61999_db
g61999_sb
g62000_da
g62000_db
g62000_sb
g62001_da
g62001_db
g62001_sb
g62002_da
g62002_db
g62002_sb
g62003_da
g62003_db
g62003_sb
g62004_sb
g62006_da
g62006_db
g62006_sb
g62007_da
g62007_db
g62007_sb
g62008_da
g62008_db
g62008_sb
g62011_da
g62011_db
g62011_sb
g62013_da
g62013_db
g62013_sb
g62015_da
g62015_db
g62015_sb
g62016_da
g62016_db
g62016_sb
g62017_da
g62017_db
g62017_sb
g62018_da
g62018_db
g62018_sb
g62021_da
g62021_db
g62021_sb
g62022_da
g62022_db
g62022_sb
g62023_da
g62023_db
g62023_sb
g62024_da
g62024_db
g62024_sb
g62026_da
g62026_db
g62026_sb
g62027_db
g62028_da
g62028_db
g62028_sb
g62029_da
g62029_db
g62029_sb
g62030_da
g62030_db
g62030_sb
g62031_da
g62031_db
g62031_sb
g62032_da
g62032_db
g62032_sb
g62033_da
g62033_db
g62033_sb
g62034_da
g62034_db
g62034_sb
g62035_da
g62035_db
g62035_sb
g62036_da
g62036_db
g62037_da
g62037_db
g62037_sb
g62038_da
g62038_db
g62038_sb
g62039_da
g62039_db
g62039_sb
g62040_da
g62040_db
g62040_sb
g62041_da
g62041_db
g62041_sb
g62042_da
g62042_db
g62042_sb
g62043_da
g62043_db
g62043_sb
g62044_da
g62044_db
g62044_sb
g62045_da
g62045_db
g62045_sb
g62046_da
g62046_db
g62048_da
g62048_db
g62048_sb
g62049_da
g62049_db
g62049_sb
g62050_da
g62050_db
g62050_sb
g62052_da
g62052_db
g62052_sb
g62053_da
g62053_db
g62053_sb
g62054_da
g62054_db
g62054_sb
g62055_da
g62055_db
g62056_da
g62056_db
g62056_sb
g62057_da
g62057_db
g62057_sb
g62058_da
g62058_db
g62058_sb
g62059_da
g62059_db
g62060_da
g62060_db
g62060_sb
g62061_da
g62061_db
g62061_sb
g62062_da
g62062_db
g62062_sb
g62063_da
g62063_db
g62063_sb
g62065_da
g62065_db
g62066_da
g62066_db
g62066_sb
g62067_da
g62067_db
g62067_sb
g62068_da
g62068_db
g62068_sb
g62069_da
g62069_db
g62069_sb
g62070_da
g62070_db
g62070_sb
g62071_da
g62071_db
g62071_sb
g62072_da
g62072_db
g62078_da
g62078_db
g62078_sb
g62079_sb
g62080_da
g62080_sb
g62081_da
g62081_db
g62081_sb
g62082_da
g62082_db
g62082_sb
g62083_da
g62083_db
g62083_sb
g62084_da
g62084_db
g62084_sb
g62085_da
g62085_db
g62085_sb
g62086_da
g62086_db
g62086_sb
g62087_da
g62087_db
g62087_sb
g62088_da
g62088_db
g62088_sb
g62089_da
g62089_db
g62089_sb
g62090_da
g62090_sb
g62091_da
g62091_db
g62091_sb
g62092_da
g62092_db
g62092_sb
g62095_da
g62095_sb
g62096_da
g62096_sb
g62097_da
g62097_sb
g62098_da
g62098_sb
g62100_da
g62100_db
g62101_da
g62101_sb
g62102_da
g62102_db
g62102_sb
g62104_da
g62104_db
g62104_sb
g62105_da
g62105_db
g62105_sb
g62106_da
g62106_db
g62106_sb
g62109_da
g62109_db
g62109_sb
g62110_da
g62110_db
g62111_da
g62111_db
g62111_sb
g62112_da
g62112_sb
g62113_da
g62113_db
g62113_sb
g62114_da
g62114_db
g62114_sb
g62116_da
g62116_db
g62117_da
g62117_sb
g62118_da
g62118_db
g62118_sb
g62119_da
g62119_db
g62120_da
g62120_sb
g62121_da
g62121_db
g62121_sb
g62122_da
g62122_db
g62122_sb
g62123_da
g62123_sb
g62124_da
g62124_sb
g62125_da
g62125_db
g62125_sb
g62126_da
g62126_sb
g62127_da
g62127_db
g62127_sb
g62128_da
g62128_db
g62128_sb
g62129_da
g62129_db
g62129_sb
g62130_da
g62130_sb
g62131_da
g62131_db
g62131_sb
g62132_da
g62132_db
g62132_sb
g62133_da
g62133_db
g62133_sb
g62134_da
g62134_db
g62134_sb
g62135_da
g62135_db
g62135_sb
g62136_da
g62136_db
g62136_sb
g62137_da
g62137_db
g62137_sb
g62138_da
g62138_sb
g62140_da
g62140_db
g62140_sb
g62219_p
g62220_p
g62221_p
g62223_p
g62254_p
g62264_p
g62266_p1
g62266_p2
g62285_p
g62312_p
g62318_p
g62326_da
g62326_db
g62326_sb
g62333_da
g62333_db
g62333_sb
g62334_da
g62334_db
g62334_sb
g62336_da
g62336_db
g62336_sb
g62339_da
g62339_db
g62339_sb
g62341_da
g62341_db
g62341_sb
g62345_da
g62345_sb
g62348_da
g62348_db
g62348_sb
g62349_da
g62349_db
g62349_sb
g62351_da
g62351_db
g62351_sb
g62352_da
g62352_db
g62352_sb
g62353_da
g62353_db
g62353_sb
g62354_da
g62354_db
g62354_sb
g62356_da
g62356_db
g62356_sb
g62357_da
g62357_db
g62357_sb
g62359_sb
g62362_db
g62362_sb
g62364_da
g62364_db
g62364_sb
g62365_da
g62365_db
g62365_sb
g62366_da
g62366_db
g62366_sb
g62367_da
g62367_db
g62367_sb
g62368_da
g62368_db
g62368_sb
g62371_da
g62371_db
g62371_sb
g62374_da
g62374_db
g62374_sb
g62375_da
g62375_db
g62375_sb
g62377_da
g62377_db
g62377_sb
g62380_da
g62380_db
g62380_sb
g62381_da
g62381_db
g62381_sb
g62383_da
g62383_db
g62383_sb
g62385_da
g62385_db
g62385_sb
g62386_da
g62386_db
g62386_sb
g62387_da
g62387_db
g62388_da
g62388_db
g62388_sb
g62389_db
g62389_sb
g62390_da
g62390_db
g62390_sb
g62391_da
g62391_db
g62391_sb
g62393_da
g62393_db
g62393_sb
g62395_da
g62395_db
g62395_sb
g62396_da
g62396_db
g62396_sb
g62398_da
g62398_db
g62398_sb
g62399_da
g62399_db
g62399_sb
g62403_da
g62403_db
g62403_sb
g62404_da
g62404_db
g62404_sb
g62406_da
g62406_db
g62406_sb
g62407_da
g62407_db
g62407_sb
g62408_da
g62408_db
g62408_sb
g62410_db
g62411_da
g62411_db
g62411_sb
g62413_da
g62413_db
g62413_sb
g62415_da
g62415_db
g62415_sb
g62419_da
g62419_sb
g62420_da
g62420_db
g62420_sb
g62422_da
g62422_db
g62422_sb
g62423_da
g62423_db
g62423_sb
g62424_da
g62424_db
g62424_sb
g62426_da
g62426_db
g62426_sb
g62427_da
g62427_db
g62427_sb
g62428_db
g62430_da
g62430_db
g62430_sb
g62431_da
g62431_db
g62431_sb
g62434_da
g62434_db
g62434_sb
g62435_da
g62435_db
g62435_sb
g62439_da
g62439_db
g62439_sb
g62440_da
g62440_db
g62440_sb
g62443_da
g62443_db
g62443_sb
g62444_da
g62444_db
g62444_sb
g62446_da
g62446_db
g62446_sb
g62447_da
g62447_db
g62447_sb
g62450_da
g62450_db
g62450_sb
g62452_da
g62452_db
g62452_sb
g62455_db
g62456_da
g62456_db
g62456_sb
g62457_da
g62457_db
g62457_sb
g62460_db
g62461_da
g62461_db
g62461_sb
g62465_da
g62465_db
g62465_sb
g62466_da
g62466_db
g62466_sb
g62467_da
g62467_db
g62467_sb
g62468_db
g62469_da
g62469_db
g62469_sb
g62470_da
g62470_db
g62470_sb
g62472_db
g62473_da
g62473_db
g62473_sb
g62475_da
g62475_db
g62475_sb
g62477_da
g62477_db
g62477_sb
g62479_da
g62479_db
g62479_sb
g62480_da
g62480_db
g62480_sb
g62481_da
g62481_db
g62482_da
g62482_db
g62482_sb
g62483_db
g62484_da
g62484_db
g62484_sb
g62485_sb
g62486_da
g62486_sb
g62487_da
g62487_db
g62487_sb
g62490_da
g62490_db
g62490_sb
g62491_da
g62491_db
g62491_sb
g62493_sb
g62494_da
g62494_db
g62494_sb
g62495_da
g62495_db
g62495_sb
g62498_da
g62498_db
g62498_sb
g62500_da
g62500_db
g62500_sb
g62502_da
g62502_db
g62502_sb
g62503_da
g62503_db
g62503_sb
g62504_da
g62504_db
g62504_sb
g62506_da
g62506_db
g62506_sb
g62509_da
g62509_db
g62509_sb
g62511_da
g62511_db
g62511_sb
g62513_da
g62513_db
g62513_sb
g62514_da
g62514_db
g62514_sb
g62517_da
g62517_db
g62517_sb
g62519_da
g62519_db
g62519_sb
g62521_da
g62521_db
g62521_sb
g62523_da
g62523_db
g62523_sb
g62527_da
g62527_db
g62527_sb
g62528_da
g62528_db
g62528_sb
g62529_da
g62529_db
g62529_sb
g62531_da
g62531_db
g62531_sb
g62532_da
g62532_db
g62532_sb
g62534_da
g62534_db
g62534_sb
g62536_da
g62536_db
g62536_sb
g62537_da
g62537_db
g62537_sb
g62538_da
g62538_sb
g62539_da
g62539_sb
g62540_da
g62540_db
g62540_sb
g62542_da
g62542_db
g62542_sb
g62544_da
g62544_db
g62544_sb
g62545_da
g62545_db
g62545_sb
g62546_da
g62546_db
g62546_sb
g62547_db
g62549_da
g62549_db
g62549_sb
g62550_da
g62550_db
g62550_sb
g62552_da
g62552_db
g62552_sb
g62554_da
g62554_db
g62554_sb
g62555_da
g62555_db
g62555_sb
g62557_da
g62557_db
g62557_sb
g62558_da
g62558_db
g62558_sb
g62559_da
g62559_db
g62559_sb
g62562_da
g62562_db
g62562_sb
g62564_da
g62564_sb
g62565_da
g62565_db
g62565_sb
g62566_da
g62566_db
g62566_sb
g62567_da
g62567_db
g62567_sb
g62568_da
g62568_db
g62568_sb
g62570_da
g62570_db
g62570_sb
g62571_da
g62571_db
g62571_sb
g62572_da
g62572_db
g62572_sb
g62574_da
g62574_db
g62574_sb
g62575_da
g62575_db
g62575_sb
g62576_da
g62576_db
g62576_sb
g62577_da
g62577_db
g62577_sb
g62580_db
g62581_da
g62581_db
g62581_sb
g62582_da
g62582_db
g62583_da
g62583_db
g62583_sb
g62585_da
g62585_db
g62585_sb
g62587_da
g62587_db
g62587_sb
g62591_da
g62591_db
g62591_sb
g62592_da
g62592_db
g62592_sb
g62593_da
g62593_db
g62593_sb
g62594_da
g62594_db
g62594_sb
g62595_p
g62596_da
g62596_db
g62596_sb
g62600_da
g62600_db
g62600_sb
g62601_sb
g62602_da
g62602_db
g62602_sb
g62604_da
g62604_db
g62604_sb
g62605_da
g62605_db
g62605_sb
g62606_da
g62606_db
g62606_sb
g62608_da
g62608_db
g62608_sb
g62610_da
g62610_db
g62610_sb
g62614_da
g62614_db
g62615_da
g62615_db
g62615_sb
g62616_da
g62616_db
g62616_sb
g62619_sb
g62622_da
g62622_db
g62622_sb
g62626_da
g62626_db
g62626_sb
g62628_da
g62628_db
g62628_sb
g62629_da
g62629_db
g62629_sb
g62630_da
g62630_db
g62630_sb
g62631_da
g62631_db
g62631_sb
g62632_da
g62632_sb
g62633_da
g62633_sb
g62634_da
g62634_db
g62634_sb
g62635_da
g62635_db
g62635_sb
g62636_da
g62636_db
g62636_sb
g62637_da
g62637_db
g62637_sb
g62638_da
g62638_db
g62638_sb
g62639_da
g62639_db
g62639_sb
g62640_da
g62640_db
g62640_sb
g62641_da
g62641_db
g62641_sb
g62643_da
g62643_db
g62643_sb
g62644_da
g62644_db
g62644_sb
g62645_da
g62645_db
g62645_sb
g62646_da
g62646_db
g62646_sb
g62647_da
g62647_db
g62647_sb
g62649_da
g62649_db
g62649_sb
g62650_da
g62650_db
g62650_sb
g62652_da
g62652_db
g62652_sb
g62653_db
g62657_da
g62657_db
g62657_sb
g62658_da
g62658_db
g62658_sb
g62659_da
g62659_db
g62659_sb
g62660_da
g62660_db
g62660_sb
g62661_da
g62661_db
g62661_sb
g62664_da
g62664_db
g62664_sb
g62666_da
g62666_db
g62666_sb
g62668_da
g62668_db
g62668_sb
g62669_da
g62669_db
g62669_sb
g62670_da
g62670_db
g62670_sb
g62672_da
g62672_db
g62672_sb
g62673_da
g62673_db
g62673_sb
g62674_da
g62674_db
g62674_sb
g62675_da
g62677_sb
g62679_da
g62679_db
g62679_sb
g62681_da
g62681_db
g62681_sb
g62683_da
g62683_db
g62683_sb
g62685_da
g62685_db
g62693_da
g62693_db
g62693_sb
g62697_db
g62698_da
g62698_db
g62698_sb
g62699_p
g62707_da
g62707_db
g62712_da
g62712_db
g62712_sb
g62714_da
g62714_db
g62714_sb
g62716_da
g62716_db
g62716_sb
g62719_da
g62719_db
g62719_sb
g62721_da
g62721_db
g62721_sb
g62723_da
g62723_db
g62723_sb
g62724_da
g62724_db
g62724_sb
g62726_da
g62726_db
g62726_sb
g62727_da
g62727_db
g62727_sb
g62729_da
g62729_db
g62729_sb
g62731_da
g62731_db
g62731_sb
g62732_da
g62732_db
g62732_sb
g62733_da
g62733_db
g62733_sb
g62735_da
g62735_db
g62735_sb
g62736_da
g62736_db
g62736_sb
g62737_da
g62737_db
g62737_sb
g62738_da
g62738_db
g62738_sb
g62739_da
g62739_db
g62739_sb
g62743_da
g62743_db
g62743_sb
g62744_da
g62744_db
g62744_sb
g62745_da
g62745_db
g62745_sb
g62746_da
g62746_db
g62746_sb
g62747_da
g62747_db
g62747_sb
g62748_da
g62748_db
g62748_sb
g62749_da
g62749_db
g62749_sb
g62750_da
g62750_db
g62750_sb
g62751_da
g62751_db
g62751_sb
g62753_da
g62753_db
g62753_sb
g62756_da
g62756_db
g62756_sb
g62757_da
g62757_db
g62757_sb
g62762_sb
g62765_da
g62765_db
g62765_sb
g62766_da
g62766_sb
g62767_da
g62767_db
g62767_sb
g62768_da
g62768_db
g62768_sb
g62769_da
g62769_db
g62769_sb
g62770_da
g62770_db
g62770_sb
g62771_da
g62771_db
g62772_da
g62772_db
g62772_sb
g62774_da
g62774_db
g62774_sb
g62775_da
g62775_db
g62775_sb
g62776_da
g62776_db
g62776_sb
g62777_da
g62777_db
g62777_sb
g62778_da
g62778_db
g62778_sb
g62782_da
g62782_db
g62782_sb
g62783_da
g62783_db
g62783_sb
g62784_da
g62784_db
g62784_sb
g62785_da
g62785_db
g62785_sb
g62786_da
g62786_db
g62786_sb
g62787_da
g62787_db
g62787_sb
g62788_da
g62788_db
g62788_sb
g62789_da
g62789_db
g62789_sb
g62791_da
g62791_db
g62791_sb
g62793_da
g62793_db
g62793_sb
g62794_da
g62794_db
g62794_sb
g62796_da
g62796_db
g62796_sb
g62797_da
g62797_db
g62797_sb
g62798_da
g62798_db
g62798_sb
g62799_da
g62799_db
g62799_sb
g62800_da
g62800_db
g62800_sb
g62802_da
g62802_db
g62802_sb
g62803_da
g62803_sb
g62804_da
g62804_db
g62804_sb
g62805_da
g62805_db
g62805_sb
g62806_da
g62806_db
g62809_da
g62809_db
g62809_sb
g62813_da
g62813_db
g62813_sb
g62814_da
g62814_db
g62814_sb
g62817_da
g62817_db
g62820_da
g62820_db
g62820_sb
g62821_da
g62821_db
g62821_sb
g62822_da
g62822_db
g62822_sb
g62824_sb
g62825_da
g62825_db
g62825_sb
g62826_da
g62826_db
g62826_sb
g62827_da
g62827_db
g62829_da
g62829_db
g62829_sb
g62830_da
g62830_db
g62830_sb
g62831_da
g62831_db
g62831_sb
g62834_da
g62834_db
g62834_sb
g62835_da
g62835_db
g62835_sb
g62836_da
g62836_db
g62836_sb
g62837_da
g62837_db
g62839_da
g62839_db
g62839_sb
g62840_da
g62840_db
g62840_sb
g62846_da
g62846_db
g62846_sb
g62847_da
g62847_db
g62847_sb
g62849_da
g62849_db
g62849_sb
g62854_da
g62854_db
g62854_sb
g62856_da
g62856_db
g62856_sb
g62857_da
g62857_db
g62857_sb
g62858_da
g62858_db
g62858_sb
g62860_da
g62860_db
g62860_sb
g62861_da
g62861_db
g62861_sb
g62862_sb
g62864_da
g62864_db
g62864_sb
g62873_p
g62874_p
g62875_p
g62876_p
g62877_p
g62879_p
g62880_p
g62881_p
g62883_da
g62883_db
g62883_sb
g62884_da
g62884_db
g62884_sb
g62885_da
g62885_db
g62885_sb
g62886_da
g62886_db
g62886_sb
g62887_da
g62887_db
g62887_sb
g62888_da
g62888_db
g62888_sb
g62889_da
g62889_db
g62889_sb
g62891_da
g62891_db
g62891_sb
g62893_da
g62893_db
g62893_sb
g62899_da
g62899_db
g62899_sb
g62900_da
g62900_db
g62900_sb
g62902_da
g62902_db
g62902_sb
g62903_da
g62903_db
g62903_sb
g62904_da
g62904_db
g62904_sb
g62905_da
g62905_db
g62905_sb
g62906_sb
g62907_da
g62907_db
g62907_sb
g62909_da
g62909_db
g62909_sb
g62911_db
g62912_da
g62912_db
g62912_sb
g62914_da
g62914_db
g62914_sb
g62915_da
g62915_db
g62915_sb
g62916_da
g62917_da
g62917_db
g62917_sb
g62918_da
g62918_db
g62918_sb
g62919_da
g62919_db
g62919_sb
g62920_da
g62920_db
g62920_sb
g62923_db
g62923_sb
g62924_da
g62924_db
g62924_sb
g62926_da
g62926_db
g62926_sb
g62929_da
g62929_db
g62929_sb
g62931_da
g62931_db
g62931_sb
g62933_da
g62933_db
g62933_sb
g62934_da
g62934_db
g62934_sb
g62935_da
g62935_db
g62935_sb
g62937_da
g62937_db
g62937_sb
g62938_da
g62938_db
g62938_sb
g62940_da
g62940_db
g62940_sb
g62941_da
g62941_db
g62941_sb
g62946_da
g62946_db
g62946_sb
g62949_da
g62949_db
g62950_da
g62950_db
g62950_sb
g62951_da
g62951_db
g62951_sb
g62953_db
g62955_da
g62955_db
g62955_sb
g62957_da
g62957_db
g62957_sb
g62959_da
g62959_db
g62959_sb
g62960_da
g62960_db
g62960_sb
g62961_da
g62961_db
g62961_sb
g62964_da
g62964_db
g62964_sb
g62969_da
g62969_db
g62969_sb
g62971_da
g62971_db
g62971_sb
g62973_da
g62973_db
g62973_sb
g62974_da
g62974_db
g62974_sb
g62976_da
g62976_db
g62976_sb
g62980_da
g62980_db
g62980_sb
g62981_da
g62981_db
g62981_sb
g62983_db
g62986_db
g62988_da
g62988_db
g62988_sb
g62989_da
g62989_db
g62989_sb
g62992_da
g62992_db
g62992_sb
g62993_da
g62993_db
g62993_sb
g63000_da
g63000_sb
g63001_da
g63001_db
g63001_sb
g63003_da
g63003_db
g63003_sb
g63008_da
g63008_db
g63008_sb
g63009_da
g63009_sb
g63010_da
g63010_db
g63010_sb
g63011_da
g63011_db
g63011_sb
g63012_da
g63012_db
g63012_sb
g63013_da
g63013_db
g63015_da
g63015_db
g63015_sb
g63016_da
g63016_db
g63016_sb
g63018_da
g63018_db
g63018_sb
g63019_da
g63019_db
g63019_sb
g63020_da
g63020_db
g63020_sb
g63024_da
g63024_db
g63027_da
g63027_db
g63027_sb
g63029_da
g63029_db
g63029_sb
g63030_da
g63030_db
g63030_sb
g63031_da
g63031_db
g63031_sb
g63034_da
g63034_db
g63034_sb
g63035_da
g63035_db
g63035_sb
g63036_da
g63036_db
g63036_sb
g63039_da
g63039_db
g63039_sb
g63040_da
g63040_db
g63040_sb
g63041_da
g63041_db
g63041_sb
g63042_da
g63042_db
g63042_sb
g63044_da
g63044_db
g63044_sb
g63045_da
g63045_db
g63045_sb
g63050_da
g63050_db
g63050_sb
g63051_da
g63051_db
g63051_sb
g63053_da
g63053_db
g63053_sb
g63054_da
g63054_db
g63054_sb
g63055_da
g63055_db
g63055_sb
g63056_da
g63056_db
g63056_sb
g63057_sb
g63058_da
g63058_sb
g63060_da
g63060_db
g63060_sb
g63063_da
g63063_db
g63063_sb
g63064_da
g63064_db
g63064_sb
g63066_da
g63066_db
g63066_sb
g63067_da
g63067_db
g63067_sb
g63069_da
g63069_db
g63069_sb
g63072_da
g63072_sb
g63073_da
g63073_db
g63073_sb
g63074_da
g63074_db
g63074_sb
g63075_da
g63075_db
g63075_sb
g63077_da
g63077_db
g63078_da
g63078_db
g63078_sb
g63079_da
g63079_db
g63079_sb
g63080_da
g63080_db
g63080_sb
g63082_da
g63082_db
g63082_sb
g63083_da
g63083_db
g63083_sb
g63086_da
g63086_db
g63086_sb
g63088_da
g63088_db
g63088_sb
g63090_da
g63090_db
g63090_sb
g63091_da
g63091_db
g63091_sb
g63093_da
g63093_db
g63093_sb
g63097_da
g63097_db
g63097_sb
g63098_da
g63098_db
g63098_sb
g63100_da
g63100_db
g63100_sb
g63101_da
g63101_db
g63101_sb
g63103_da
g63103_db
g63103_sb
g63105_da
g63105_db
g63105_sb
g63106_da
g63106_db
g63106_sb
g63108_da
g63108_db
g63108_sb
g63109_da
g63109_db
g63109_sb
g63110_da
g63110_db
g63110_sb
g63113_da
g63113_db
g63113_sb
g63114_da
g63114_db
g63114_sb
g63115_da
g63115_db
g63115_sb
g63116_da
g63116_db
g63116_sb
g63117_da
g63117_db
g63117_sb
g63118_da
g63118_db
g63118_sb
g63119_da
g63119_db
g63119_sb
g63122_da
g63122_sb
g63123_da
g63123_db
g63123_sb
g63125_da
g63125_db
g63125_sb
g63127_da
g63127_db
g63127_sb
g63128_da
g63128_db
g63128_sb
g63130_da
g63130_db
g63130_sb
g63132_da
g63132_db
g63132_sb
g63133_da
g63133_db
g63134_da
g63134_db
g63134_sb
g63135_da
g63135_db
g63135_sb
g63137_da
g63137_db
g63137_sb
g63138_da
g63138_db
g63138_sb
g63142_da
g63142_db
g63142_sb
g63145_da
g63145_db
g63145_sb
g63146_da
g63146_db
g63146_sb
g63148_da
g63148_db
g63148_sb
g63149_da
g63149_db
g63149_sb
g63150_da
g63150_db
g63150_sb
g63151_da
g63151_db
g63151_sb
g63154_sb
g63158_db
g63158_sb
g63163_da
g63163_db
g63163_sb
g63166_da
g63166_db
g63166_sb
g63168_da
g63168_db
g63168_sb
g63169_da
g63169_db
g63169_sb
g63172_da
g63172_db
g63172_sb
g63173_da
g63173_db
g63173_sb
g63175_da
g63175_db
g63175_sb
g63179_da
g63179_db
g63179_sb
g63180_da
g63180_db
g63180_sb
g63181_da
g63181_db
g63181_sb
g63182_da
g63182_db
g63182_sb
g63183_da
g63183_sb
g63184_db
g63184_sb
g63186_da
g63186_db
g63186_sb
g63187_da
g63187_db
g63187_sb
g63188_da
g63188_db
g63188_sb
g63189_da
g63189_db
g63189_sb
g63190_da
g63190_db
g63190_sb
g63193_da
g63193_db
g63193_sb
g63194_da
g63194_db
g63194_sb
g63195_da
g63195_db
g63195_sb
g63196_da
g63196_db
g63196_sb
g63197_da
g63197_db
g63197_sb
g63198_da
g63198_db
g63198_sb
g63199_da
g63199_db
g63199_sb
g63200_p
g63201_p
g63202_da
g63202_db
g63202_sb
g63203_da
g63203_db
g63203_sb
g63204_da
g63204_db
g63204_sb
g63207_p
g63209_p
g63216_p
g63217_p
g63253_p
g63256_p
g63259_p
g63263_p
g63271_p
g63291_p
g63292_p
g63293_p
g63340_p
g63348_p
g63364_p
g63378_da
g63378_db
g63378_sb
g63392_da
g63392_db
g63392_sb
g63397_da
g63397_db
g63397_sb
g63409_p
g63422_p
g63423_p
g63424_p
g63426_p
g63429_p
g63430_p
g63431_da
g63431_db
g63431_sb
g63432_da
g63432_db
g63432_sb
g63433_da
g63433_db
g63433_sb
g63434_da
g63434_db
g63434_sb
g63435_da
g63435_db
g63435_sb
g63436_da
g63436_db
g63436_sb
g63437_da
g63437_db
g63437_sb
g63438_da
g63438_db
g63438_sb
g63525_p
g63539_p
g63542_p
g63546_p
g63547_da
g63547_db
g63547_sb
g63550_da
g63550_db
g63550_sb
g63551_da
g63551_db
g63551_sb
g63552_da
g63552_db
g63552_sb
g63553_da
g63553_db
g63553_sb
g63554_da
g63554_db
g63554_sb
g63555_da
g63555_db
g63555_sb
g63556_da
g63556_db
g63556_sb
g63557_da
g63557_db
g63557_sb
g63559_da
g63559_db
g63559_sb
g63560_da
g63560_db
g63560_sb
g63561_da
g63561_db
g63561_sb
g63562_da
g63562_db
g63562_sb
g63564_sb
g63567_da
g63567_db
g63567_sb
g63568_da
g63568_db
g63568_sb
g63569_da
g63569_db
g63569_sb
g63570_da
g63570_db
g63570_sb
g63571_da
g63571_db
g63571_sb
g63572_da
g63572_db
g63572_sb
g63573_da
g63573_db
g63573_sb
g63574_da
g63574_db
g63574_sb
g63576_da
g63576_db
g63576_sb
g63577_da
g63577_db
g63577_sb
g63578_p
g63579_p
g63580_p
g63581_p
g63582_da
g63582_db
g63582_sb
g63583_da
g63583_db
g63583_sb
g63585_da
g63587_db
g63588_da
g63588_db
g63588_sb
g63589_da
g63589_db
g63589_sb
g63590_da
g63590_db
g63590_sb
g63591_da
g63591_db
g63591_sb
g63592_da
g63592_db
g63592_sb
g63593_da
g63593_db
g63593_sb
g63594_da
g63594_db
g63594_sb
g63595_da
g63595_db
g63595_sb
g63596_da
g63596_db
g63596_sb
g63597_da
g63597_db
g63597_sb
g63598_da
g63598_db
g63598_sb
g63599_da
g63599_db
g63599_sb
g63600_da
g63600_db
g63600_sb
g63601_da
g63601_db
g63601_sb
g63602_da
g63602_db
g63602_sb
g63603_da
g63603_db
g63603_sb
g63604_da
g63604_db
g63604_sb
g63605_da
g63605_db
g63605_sb
g63606_da
g63606_db
g63606_sb
g63607_da
g63607_db
g63607_sb
g63608_da
g63608_db
g63608_sb
g63609_da
g63609_db
g63609_sb
g63610_da
g63610_db
g63610_sb
g63611_da
g63611_db
g63611_sb
g63612_da
g63612_db
g63612_sb
g63613_da
g63613_db
g63613_sb
g63614_da
g63614_db
g63614_sb
g63615_da
g63615_db
g63615_sb
g63616_da
g63616_db
g63616_sb
g63617_da
g63617_db
g63617_sb
g63618_da
g63618_db
g63618_sb
g63619_da
g63619_db
g63619_sb
g63620_da
g63620_db
g63620_sb
g63621_da
g63621_db
g63621_sb
g63891_p
g63892_p
g63901_p
g63902_p
g63916_p
g63922_p
g63939_p
g63943_AP
g63943_BP
g63943_p
g64078_da
g64078_sb
g64079_da
g64079_db
g64079_sb
g64081_da
g64081_db
g64081_sb
g64082_da
g64082_db
g64082_sb
g64084_da
g64084_db
g64084_sb
g64090_da
g64090_db
g64090_sb
g64094_da
g64094_db
g64094_sb
g64095_da
g64095_db
g64095_sb
g64097_da
g64097_db
g64097_sb
g64099_da
g64099_db
g64099_sb
g64102_da
g64102_db
g64102_sb
g64103_da
g64103_db
g64103_sb
g64106_da
g64106_db
g64106_sb
g64107_da
g64107_db
g64107_sb
g64108_da
g64108_db
g64108_sb
g64109_da
g64109_db
g64109_sb
g64110_da
g64110_db
g64110_sb
g64111_da
g64111_db
g64111_sb
g64113_da
g64113_db
g64113_sb
g64114_da
g64114_db
g64114_sb
g64115_da
g64115_db
g64115_sb
g64117_da
g64117_db
g64117_sb
g64119_da
g64119_db
g64122_da
g64122_db
g64124_p
g64125_da
g64125_db
g64125_sb
g64126_da
g64126_db
g64126_sb
g64127_da
g64127_db
g64127_sb
g64130_da
g64130_db
g64130_sb
g64131_da
g64131_db
g64131_sb
g64132_da
g64132_db
g64132_sb
g64133_da
g64133_db
g64133_sb
g64138_da
g64138_db
g64138_sb
g64139_da
g64139_db
g64139_sb
g64140_da
g64140_db
g64140_sb
g64141_da
g64141_db
g64141_sb
g64142_da
g64142_db
g64142_sb
g64143_da
g64143_db
g64143_sb
g64145_da
g64145_db
g64145_sb
g64146_da
g64146_db
g64146_sb
g64148_da
g64148_db
g64149_da
g64149_db
g64149_sb
g64152_da
g64152_db
g64152_sb
g64153_da
g64153_db
g64153_sb
g64156_da
g64156_db
g64156_sb
g64157_da
g64157_db
g64158_da
g64158_db
g64158_sb
g64162_da
g64162_db
g64163_da
g64163_db
g64163_sb
g64165_da
g64165_db
g64165_sb
g64168_da
g64168_db
g64168_sb
g64169_da
g64169_db
g64169_sb
g64170_da
g64170_db
g64170_sb
g64171_da
g64171_db
g64171_sb
g64172_da
g64172_db
g64172_sb
g64175_da
g64175_db
g64175_sb
g64176_da
g64176_db
g64177_da
g64177_db
g64177_sb
g64178_da
g64178_db
g64178_sb
g64179_da
g64179_db
g64179_sb
g64182_da
g64182_db
g64182_sb
g64184_da
g64184_db
g64185_da
g64185_db
g64185_sb
g64187_da
g64187_db
g64187_sb
g64188_da
g64188_db
g64188_sb
g64189_da
g64189_db
g64189_sb
g64190_da
g64190_db
g64190_sb
g64192_da
g64192_db
g64192_sb
g64194_p
g64196_da
g64196_db
g64196_sb
g64200_da
g64200_db
g64200_sb
g64201_da
g64201_db
g64201_sb
g64202_da
g64202_db
g64202_sb
g64204_da
g64204_db
g64204_sb
g64208_da
g64208_db
g64208_sb
g64209_da
g64209_db
g64209_sb
g64210_da
g64210_db
g64210_sb
g64211_da
g64211_db
g64211_sb
g64213_da
g64213_db
g64213_sb
g64214_da
g64214_db
g64214_sb
g64215_da
g64215_db
g64215_sb
g64216_da
g64216_db
g64216_sb
g64217_db
g64217_sb
g64219_da
g64219_db
g64219_sb
g64222_da
g64222_db
g64222_sb
g64223_da
g64223_sb
g64224_da
g64224_db
g64224_sb
g64225_da
g64225_db
g64225_sb
g64226_da
g64226_db
g64226_sb
g64227_da
g64227_db
g64227_sb
g64231_da
g64231_db
g64231_sb
g64232_da
g64232_db
g64232_sb
g64235_da
g64235_db
g64237_da
g64237_db
g64237_sb
g64239_da
g64239_db
g64239_sb
g64243_da
g64243_db
g64243_sb
g64244_da
g64244_db
g64244_sb
g64245_da
g64245_db
g64245_sb
g64246_da
g64246_db
g64246_sb
g64251_da
g64251_db
g64251_sb
g64252_da
g64252_db
g64252_sb
g64255_da
g64255_db
g64255_sb
g64256_da
g64256_db
g64256_sb
g64259_da
g64259_db
g64259_sb
g64264_da
g64264_db
g64264_sb
g64267_da
g64267_db
g64267_sb
g64268_da
g64268_db
g64268_sb
g64269_da
g64269_db
g64269_sb
g64272_da
g64272_db
g64272_sb
g64273_da
g64273_db
g64276_da
g64276_db
g64276_sb
g64278_da
g64278_db
g64278_sb
g64280_da
g64280_db
g64280_sb
g64282_da
g64282_db
g64282_sb
g64284_da
g64284_db
g64284_sb
g64286_da
g64286_db
g64286_sb
g64288_da
g64288_db
g64288_sb
g64289_da
g64289_db
g64289_sb
g64290_da
g64290_db
g64290_sb
g64291_da
g64291_db
g64291_sb
g64294_da
g64294_db
g64294_sb
g64295_da
g64295_db
g64295_sb
g64296_db
g64297_da
g64297_db
g64297_sb
g64298_da
g64298_db
g64298_sb
g64300_da
g64300_db
g64300_sb
g64301_da
g64301_db
g64301_sb
g64303_da
g64303_db
g64303_sb
g64305_da
g64305_db
g64305_sb
g64309_da
g64309_db
g64309_sb
g64310_da
g64310_db
g64310_sb
g64311_da
g64311_db
g64311_sb
g64312_da
g64312_db
g64312_sb
g64313_da
g64313_db
g64315_da
g64315_db
g64315_sb
g64316_da
g64316_db
g64316_sb
g64320_da
g64320_db
g64320_sb
g64322_da
g64322_db
g64322_sb
g64323_da
g64323_db
g64323_sb
g64324_da
g64324_db
g64324_sb
g64325_da
g64325_db
g64325_sb
g64326_db
g64326_sb
g64327_da
g64327_db
g64327_sb
g64329_da
g64329_db
g64329_sb
g64331_da
g64331_db
g64331_sb
g64332_da
g64332_db
g64332_sb
g64333_da
g64333_db
g64333_sb
g64339_da
g64339_db
g64339_sb
g64343_da
g64343_db
g64343_sb
g64344_da
g64344_db
g64344_sb
g64345_da
g64345_db
g64345_sb
g64346_da
g64346_db
g64346_sb
g64348_da
g64348_db
g64348_sb
g64349_da
g64349_db
g64349_sb
g64351_da
g64351_db
g64351_sb
g64354_da
g64354_db
g64354_sb
g64355_da
g64355_db
g64355_sb
g64356_da
g64356_db
g64356_sb
g64358_da
g64358_db
g64358_sb
g64359_da
g64359_db
g64359_sb
g64360_da
g64360_db
g64360_sb
g64362_da
g64362_db
g64362_sb
g64363_da
g64363_db
g64363_sb
g64365_db
g64367_da
g64367_db
g64367_sb
g64368_p
g64369_p
g64370_p
g64375_p
g64376_p
g64377_p
g64378_p
g64379_p
g64380_p
g64383_p
g64384_p
g64454_p
g64461_p
g64465_p
g64466_p
g64577_p
g64578_p
g64581_p
g64582_p
g64585_p
g64587_p
g64595_p
g64596_p
g64610_p
g64630_AP
g64630_BP
g64630_p
g64631_p
g64633_p
g64639_p
g64643_p
g64646_p
g64671_p
g64678_p
g64687_p
g64697_p
g64700_p
g64701_p
g64702_p
g64704_p
g64705_p
g64712_p
g64727_p
g64736_p
g64740_p
g64746_p
g64747_p
g64748_da
g64748_db
g64748_sb
g64749_da
g64749_db
g64752_da
g64752_db
g64752_sb
g64754_da
g64754_db
g64754_sb
g64756_da
g64756_db
g64756_sb
g64758_da
g64758_db
g64758_sb
g64760_da
g64760_db
g64760_sb
g64763_da
g64763_db
g64763_sb
g64764_da
g64764_db
g64764_sb
g64765_da
g64765_db
g64767_da
g64767_db
g64767_sb
g64768_da
g64768_db
g64768_sb
g64769_da
g64769_db
g64769_sb
g64770_da
g64770_db
g64770_sb
g64772_da
g64772_db
g64772_sb
g64773_da
g64773_db
g64773_sb
g64775_da
g64775_db
g64775_sb
g64776_db
g64777_da
g64777_db
g64777_sb
g64780_da
g64780_db
g64780_sb
g64781_da
g64781_db
g64781_sb
g64784_da
g64784_db
g64784_sb
g64786_da
g64786_db
g64786_sb
g64788_da
g64788_db
g64788_sb
g64790_da
g64790_db
g64790_sb
g64791_da
g64791_db
g64791_sb
g64793_da
g64793_db
g64793_sb
g64797_da
g64797_db
g64797_sb
g64799_da
g64799_db
g64799_sb
g64800_sb
g64808_da
g64808_db
g64808_sb
g64809_da
g64809_db
g64809_sb
g64811_da
g64811_db
g64811_sb
g64813_da
g64813_db
g64813_sb
g64814_da
g64814_db
g64814_sb
g64816_da
g64816_db
g64816_sb
g64818_da
g64818_db
g64818_sb
g64821_da
g64821_db
g64821_sb
g64826_da
g64826_sb
g64827_da
g64827_db
g64827_sb
g64829_da
g64829_db
g64829_sb
g64833_da
g64833_db
g64833_sb
g64834_da
g64834_db
g64834_sb
g64835_da
g64835_db
g64835_sb
g64836_da
g64836_db
g64836_sb
g64839_da
g64839_sb
g64840_da
g64842_da
g64842_db
g64842_sb
g64844_da
g64844_db
g64844_sb
g64845_da
g64845_db
g64845_sb
g64847_da
g64847_db
g64847_sb
g64850_da
g64850_db
g64850_sb
g64851_da
g64851_db
g64851_sb
g64852_da
g64852_db
g64852_sb
g64854_da
g64854_db
g64854_sb
g64855_da
g64855_db
g64855_sb
g64856_da
g64856_db
g64856_sb
g64857_da
g64857_db
g64857_sb
g64859_da
g64859_db
g64859_sb
g64861_sb
g64863_da
g64863_db
g64863_sb
g64864_da
g64864_db
g64864_sb
g64866_da
g64866_db
g64866_sb
g64867_da
g64867_db
g64867_sb
g64872_da
g64872_db
g64872_sb
g64874_da
g64874_db
g64875_da
g64875_db
g64875_sb
g64876_da
g64876_db
g64876_sb
g64877_da
g64877_db
g64877_sb
g64880_da
g64880_db
g64880_sb
g64881_da
g64881_db
g64881_sb
g64883_da
g64883_db
g64883_sb
g64884_da
g64884_sb
g64885_da
g64885_db
g64885_sb
g64886_da
g64886_db
g64886_sb
g64887_da
g64887_db
g64887_sb
g64888_da
g64888_db
g64889_da
g64889_db
g64889_sb
g64890_da
g64890_db
g64890_sb
g64891_da
g64891_db
g64891_sb
g64893_da
g64893_db
g64893_sb
g64894_da
g64894_db
g64894_sb
g64896_da
g64896_db
g64896_sb
g64897_da
g64897_db
g64897_sb
g64898_da
g64898_db
g64898_sb
g64899_da
g64899_db
g64899_sb
g64904_da
g64904_db
g64904_sb
g64905_da
g64905_db
g64905_sb
g64906_sb
g64907_sb
g64908_da
g64908_sb
g64910_da
g64910_db
g64910_sb
g64911_da
g64911_db
g64911_sb
g64919_da
g64919_db
g64919_sb
g64921_da
g64921_db
g64921_sb
g64925_da
g64925_db
g64925_sb
g64927_da
g64927_db
g64927_sb
g64928_db
g64929_db
g64930_da
g64930_db
g64930_sb
g64931_da
g64931_db
g64931_sb
g64933_da
g64933_db
g64933_sb
g64934_da
g64934_db
g64934_sb
g64936_da
g64936_db
g64936_sb
g64937_da
g64937_db
g64937_sb
g64938_da
g64938_db
g64938_sb
g64939_da
g64939_sb
g64940_da
g64940_db
g64940_sb
g64941_da
g64941_db
g64941_sb
g64943_da
g64943_db
g64943_sb
g64944_da
g64944_db
g64945_da
g64945_db
g64945_sb
g64947_da
g64947_db
g64947_sb
g64948_da
g64948_sb
g64949_da
g64949_db
g64949_sb
g64950_da
g64950_db
g64950_sb
g64951_da
g64951_db
g64951_sb
g64952_da
g64952_db
g64952_sb
g64954_da
g64954_db
g64954_sb
g64957_da
g64957_db
g64957_sb
g64958_da
g64958_db
g64958_sb
g64959_da
g64959_db
g64959_sb
g64962_da
g64962_db
g64962_sb
g64965_da
g64965_db
g64965_sb
g64966_da
g64966_db
g64967_da
g64967_db
g64967_sb
g64969_da
g64969_db
g64969_sb
g64971_da
g64971_db
g64971_sb
g64974_da
g64974_db
g64976_da
g64976_db
g64976_sb
g64979_da
g64979_db
g64979_sb
g64980_da
g64980_db
g64980_sb
g64984_da
g64984_db
g64984_sb
g64986_da
g64986_db
g64986_sb
g64987_da
g64987_db
g64987_sb
g64989_da
g64989_sb
g64992_da
g64992_db
g64992_sb
g64993_db
g64994_da
g64994_db
g64997_da
g64997_db
g64997_sb
g64998_da
g64998_db
g64998_sb
g64999_da
g64999_db
g64999_sb
g65000_da
g65000_db
g65000_sb
g65002_da
g65002_db
g65002_sb
g65003_da
g65003_db
g65003_sb
g65004_db
g65005_da
g65005_db
g65005_sb
g65006_da
g65006_db
g65006_sb
g65007_da
g65007_db
g65007_sb
g65009_da
g65009_db
g65011_da
g65011_db
g65011_sb
g65012_da
g65012_db
g65012_sb
g65013_da
g65013_db
g65013_sb
g65015_db
g65016_da
g65016_db
g65016_sb
g65019_da
g65019_db
g65019_sb
g65020_da
g65020_db
g65020_sb
g65021_db
g65022_db
g65022_sb
g65023_da
g65023_db
g65023_sb
g65024_da
g65024_db
g65024_sb
g65025_da
g65025_db
g65025_sb
g65026_da
g65026_db
g65026_sb
g65027_da
g65027_db
g65027_sb
g65029_da
g65029_db
g65029_sb
g65030_da
g65030_db
g65030_sb
g65032_da
g65032_db
g65032_sb
g65033_da
g65033_db
g65033_sb
g65035_da
g65035_db
g65035_sb
g65037_da
g65037_db
g65037_sb
g65038_da
g65038_db
g65038_sb
g65039_da
g65039_db
g65039_sb
g65040_da
g65040_db
g65040_sb
g65041_da
g65041_db
g65041_sb
g65042_da
g65042_db
g65042_sb
g65044_da
g65044_db
g65044_sb
g65045_da
g65045_db
g65045_sb
g65047_da
g65047_db
g65047_sb
g65053_da
g65053_db
g65053_sb
g65054_da
g65054_db
g65054_sb
g65055_da
g65055_db
g65055_sb
g65056_da
g65056_db
g65056_sb
g65058_da
g65058_db
g65058_sb
g65059_da
g65059_sb
g65060_da
g65060_db
g65060_sb
g65064_da
g65064_db
g65064_sb
g65066_da
g65066_db
g65066_sb
g65067_da
g65067_db
g65067_sb
g65069_da
g65069_db
g65069_sb
g65077_da
g65077_db
g65077_sb
g65078_da
g65078_db
g65078_sb
g65079_da
g65079_db
g65079_sb
g65081_da
g65081_db
g65081_sb
g65082_da
g65082_sb
g65083_da
g65083_db
g65083_sb
g65084_da
g65084_db
g65084_sb
g65085_da
g65085_db
g65085_sb
g65086_da
g65086_db
g65086_sb
g65087_da
g65087_db
g65091_da
g65091_db
g65091_sb
g65092_da
g65092_sb
g65093_da
g65093_db
g65093_sb
g65094_da
g65094_db
g65094_sb
g65095_da
g65095_db
g65095_sb
g65096_da
g65096_db
g65096_sb
g65097_da
g65097_db
g65097_sb
g65210_da
g65210_db
g65210_sb
g65211_da
g65211_db
g65211_sb
g65212_da
g65212_db
g65213_da
g65213_db
g65213_sb
g65214_da
g65214_db
g65214_sb
g65215_da
g65216_da
g65216_db
g65216_sb
g65217_da
g65217_db
g65217_sb
g65221_da
g65221_db
g65221_sb
g65222_da
g65222_db
g65222_sb
g65223_da
g65223_db
g65223_sb
g65224_da
g65224_db
g65224_sb
g65225_da
g65225_sb
g65226_da
g65226_db
g65226_sb
g65228_da
g65228_db
g65228_sb
g65230_da
g65230_db
g65230_sb
g65232_da
g65232_db
g65232_sb
g65233_da
g65233_db
g65233_sb
g65234_da
g65234_sb
g65235_da
g65235_db
g65235_sb
g65236_da
g65236_db
g65236_sb
g65237_da
g65237_db
g65237_sb
g65238_da
g65238_db
g65238_sb
g65240_da
g65240_db
g65240_sb
g65241_da
g65241_db
g65241_sb
g65242_da
g65242_db
g65242_sb
g65243_da
g65243_db
g65243_sb
g65244_da
g65244_db
g65244_sb
g65245_da
g65245_db
g65245_sb
g65246_da
g65246_db
g65246_sb
g65247_da
g65247_db
g65247_sb
g65248_da
g65248_db
g65248_sb
g65249_da
g65249_db
g65249_sb
g65250_da
g65250_db
g65250_sb
g65251_da
g65251_db
g65251_sb
g65252_da
g65252_db
g65252_sb
g65254_p
g65255_p
g65256_da
g65256_db
g65257_p
g65258_p
g65259_p
g65260_p
g65262_da
g65262_db
g65262_sb
g65263_p
g65264_p
g65265_p
g65266_p
g65267_p
g65268_da
g65268_db
g65268_sb
g65270_da
g65270_db
g65270_sb
g65271_da
g65271_db
g65271_sb
g65272_da
g65272_db
g65272_sb
g65274_da
g65274_db
g65274_sb
g65277_da
g65277_db
g65277_sb
g65280_da
g65280_db
g65280_sb
g65281_da
g65281_db
g65281_sb
g65282_da
g65282_db
g65282_sb
g65283_da
g65283_db
g65283_sb
g65284_da
g65284_db
g65284_sb
g65285_da
g65285_db
g65285_sb
g65286_da
g65286_db
g65286_sb
g65288_da
g65288_db
g65288_sb
g65289_da
g65289_db
g65289_sb
g65291_da
g65291_db
g65291_sb
g65293_da
g65293_db
g65293_sb
g65295_da
g65295_db
g65295_sb
g65297_da
g65297_db
g65297_sb
g65299_da
g65299_db
g65299_sb
g65300_da
g65300_db
g65300_sb
g65301_da
g65302_da
g65302_db
g65302_sb
g65303_da
g65303_db
g65303_sb
g65304_da
g65304_db
g65304_sb
g65305_sb
g65306_da
g65306_db
g65306_sb
g65307_da
g65307_db
g65307_sb
g65310_da
g65310_db
g65310_sb
g65314_da
g65314_sb
g65316_da
g65316_db
g65316_sb
g65317_da
g65317_db
g65317_sb
g65318_da
g65318_db
g65318_sb
g65319_da
g65319_db
g65319_sb
g65323_da
g65323_db
g65323_sb
g65325_da
g65325_db
g65327_da
g65327_db
g65327_sb
g65328_da
g65328_db
g65328_sb
g65329_sb
g65331_da
g65331_db
g65331_sb
g65332_da
g65332_db
g65332_sb
g65334_da
g65334_db
g65335_da
g65336_da
g65336_db
g65336_sb
g65337_da
g65337_db
g65337_sb
g65338_da
g65338_db
g65338_sb
g65339_da
g65339_db
g65339_sb
g65341_da
g65341_db
g65341_sb
g65342_da
g65342_db
g65342_sb
g65345_da
g65345_db
g65345_sb
g65346_da
g65346_db
g65346_sb
g65348_da
g65348_db
g65348_sb
g65349_da
g65349_db
g65349_sb
g65350_da
g65350_db
g65350_sb
g65351_sb
g65354_da
g65354_db
g65354_sb
g65356_da
g65356_db
g65356_sb
g65357_sb
g65358_da
g65358_db
g65358_sb
g65359_da
g65359_db
g65359_sb
g65360_da
g65360_db
g65360_sb
g65364_da
g65364_db
g65364_sb
g65368_da
g65368_sb
g65369_db
g65369_sb
g65371_da
g65371_db
g65371_sb
g65372_da
g65372_db
g65372_sb
g65373_da
g65373_db
g65373_sb
g65376_da
g65376_db
g65376_sb
g65377_da
g65377_db
g65377_sb
g65380_da
g65380_db
g65380_sb
g65381_db
g65386_da
g65386_db
g65386_sb
g65387_da
g65387_db
g65387_sb
g65388_da
g65388_db
g65388_sb
g65389_da
g65389_db
g65389_sb
g65390_da
g65390_db
g65390_sb
g65391_da
g65391_db
g65391_sb
g65393_da
g65393_db
g65393_sb
g65394_da
g65394_db
g65394_sb
g65399_da
g65399_db
g65399_sb
g65403_da
g65403_db
g65403_sb
g65404_da
g65404_db
g65404_sb
g65406_da
g65406_db
g65406_sb
g65408_da
g65408_db
g65408_sb
g65409_da
g65409_db
g65409_sb
g65411_da
g65411_db
g65411_sb
g65416_da
g65416_db
g65416_sb
g65418_da
g65418_db
g65418_sb
g65420_da
g65420_db
g65420_sb
g65423_da
g65423_db
g65423_sb
g65425_da
g65425_db
g65425_sb
g65426_da
g65426_db
g65426_sb
g65427_da
g65427_db
g65427_sb
g65428_da
g65428_db
g65428_sb
g65429_da
g65429_db
g65429_sb
g65431_da
g65431_db
g65431_sb
g65435_da
g65435_db
g65435_sb
g65436_p
g65437_p
g65439_p
g65486_p
g65488_p
g65489_p
g65490_p
g65491_p
g65495_p
g65496_p
g65497_p
g65498_p
g65511_p
g65513_p
g65514_p
g65515_p
g65517_p
g65518_p
g65530_p
g65533_p
g65543_p
g65549_p
g65550_p
g65557_p
g65559_p
g65562_p
g65567_p
g65568_p
g65569_p
g65570_p
g65571_p
g65572_p1
g65572_p2
g65583_p
g65588_p
g65590_p
g65595_p
g65614_p
g65617_p
g65626_p
g65674_da
g65674_db
g65674_sb
g65675_da
g65675_db
g65675_sb
g65677_da
g65677_db
g65677_sb
g65678_da
g65678_db
g65678_sb
g65679_da
g65679_db
g65679_sb
g65680_da
g65680_db
g65680_sb
g65681_da
g65681_db
g65681_sb
g65684_da
g65684_db
g65684_sb
g65685_da
g65685_db
g65685_sb
g65686_da
g65686_db
g65686_sb
g65687_da
g65687_db
g65687_sb
g65688_da
g65688_db
g65688_sb
g65689_da
g65689_db
g65689_sb
g65691_da
g65691_db
g65691_sb
g65692_da
g65692_db
g65692_sb
g65693_da
g65693_db
g65693_sb
g65694_da
g65694_db
g65694_sb
g65696_da
g65696_db
g65696_sb
g65697_da
g65697_db
g65697_sb
g65699_da
g65699_db
g65699_sb
g65700_da
g65700_db
g65700_sb
g65701_da
g65701_db
g65701_sb
g65702_da
g65702_db
g65702_sb
g65703_da
g65703_db
g65703_sb
g65704_da
g65704_db
g65704_sb
g65705_da
g65705_db
g65705_sb
g65709_da
g65709_db
g65709_sb
g65711_da
g65711_db
g65711_sb
g65712_da
g65712_db
g65712_sb
g65713_da
g65713_db
g65713_sb
g65714_da
g65714_db
g65714_sb
g65715_da
g65715_db
g65715_sb
g65716_da
g65716_db
g65716_sb
g65717_da
g65717_db
g65717_sb
g65718_da
g65718_db
g65718_sb
g65719_da
g65719_db
g65719_sb
g65720_da
g65720_db
g65720_sb
g65721_da
g65721_db
g65721_sb
g65723_da
g65723_db
g65723_sb
g65724_da
g65724_db
g65724_sb
g65725_da
g65725_db
g65725_sb
g65726_da
g65726_db
g65726_sb
g65727_da
g65727_db
g65727_sb
g65728_da
g65728_db
g65728_sb
g65729_p
g65730_da
g65730_db
g65730_sb
g65732_da
g65732_db
g65732_sb
g65733_da
g65733_db
g65733_sb
g65734_da
g65734_db
g65734_sb
g65736_da
g65736_db
g65736_sb
g65737_da
g65737_db
g65737_sb
g65740_da
g65740_db
g65740_sb
g65741_da
g65741_db
g65741_sb
g65743_da
g65743_db
g65743_sb
g65744_da
g65744_db
g65744_sb
g65745_da
g65745_db
g65745_sb
g65746_da
g65746_db
g65746_sb
g65748_da
g65748_db
g65748_sb
g65749_da
g65749_db
g65749_sb
g65752_da
g65752_db
g65752_sb
g65753_da
g65753_db
g65753_sb
g65754_da
g65754_db
g65754_sb
g65756_da
g65756_db
g65756_sb
g65757_da
g65757_db
g65757_sb
g65759_da
g65759_db
g65759_sb
g65760_da
g65760_db
g65760_sb
g65761_da
g65761_db
g65761_sb
g65762_da
g65762_db
g65762_sb
g65763_da
g65763_db
g65763_sb
g65764_da
g65764_db
g65764_sb
g65765_da
g65765_db
g65765_sb
g65766_da
g65766_db
g65766_sb
g65767_da
g65767_db
g65767_sb
g65768_da
g65768_db
g65768_sb
g65769_da
g65769_db
g65769_sb
g65770_da
g65770_db
g65770_sb
g65772_da
g65772_db
g65772_sb
g65774_da
g65774_db
g65774_sb
g65776_da
g65776_db
g65776_sb
g65777_da
g65777_db
g65777_sb
g65778_da
g65778_db
g65778_sb
g65779_da
g65779_db
g65779_sb
g65780_da
g65780_db
g65780_sb
g65781_da
g65781_db
g65781_sb
g65782_da
g65782_db
g65782_sb
g65783_da
g65783_db
g65783_sb
g65784_da
g65784_db
g65784_sb
g65785_da
g65785_db
g65785_sb
g65787_da
g65787_db
g65787_sb
g65788_da
g65788_db
g65788_sb
g65790_da
g65790_db
g65790_sb
g65791_da
g65791_db
g65791_sb
g65792_da
g65792_db
g65792_sb
g65793_da
g65793_db
g65793_sb
g65794_da
g65794_db
g65794_sb
g65795_da
g65795_db
g65795_sb
g65796_da
g65796_db
g65796_sb
g65799_da
g65799_db
g65799_sb
g65800_da
g65800_db
g65800_sb
g65801_p
g65802_da
g65802_db
g65802_sb
g65803_da
g65803_db
g65803_sb
g65805_da
g65805_db
g65805_sb
g65807_da
g65807_db
g65807_sb
g65809_da
g65809_db
g65809_sb
g65810_da
g65810_db
g65810_sb
g65811_da
g65811_db
g65811_sb
g65812_da
g65812_db
g65812_sb
g65813_da
g65813_db
g65813_sb
g65814_da
g65814_db
g65814_sb
g65816_da
g65816_db
g65816_sb
g65817_da
g65817_db
g65817_sb
g65819_da
g65819_db
g65819_sb
g65822_da
g65822_db
g65822_sb
g65823_db
g65824_da
g65824_db
g65824_sb
g65825_da
g65825_db
g65825_sb
g65826_da
g65826_db
g65826_sb
g65827_da
g65827_db
g65827_sb
g65828_da
g65828_db
g65828_sb
g65829_da
g65829_db
g65829_sb
g65830_da
g65830_db
g65830_sb
g65831_da
g65831_db
g65831_sb
g65832_da
g65832_db
g65832_sb
g65833_da
g65833_db
g65833_sb
g65834_da
g65834_db
g65834_sb
g65835_da
g65835_db
g65835_sb
g65837_da
g65837_db
g65837_sb
g65838_da
g65838_db
g65838_sb
g65840_da
g65840_db
g65840_sb
g65843_da
g65843_db
g65843_sb
g65844_da
g65844_db
g65844_sb
g65846_da
g65846_db
g65846_sb
g65847_da
g65847_db
g65847_sb
g65849_da
g65849_db
g65849_sb
g65850_da
g65850_db
g65850_sb
g65852_da
g65852_db
g65852_sb
g65853_da
g65853_db
g65853_sb
g65855_da
g65855_db
g65855_sb
g65856_da
g65856_db
g65856_sb
g65857_da
g65857_db
g65857_sb
g65858_da
g65858_db
g65858_sb
g65860_da
g65860_db
g65860_sb
g65861_da
g65861_db
g65861_sb
g65863_da
g65863_db
g65863_sb
g65865_da
g65865_db
g65865_sb
g65866_da
g65866_db
g65866_sb
g65867_da
g65867_db
g65867_sb
g65870_da
g65870_db
g65870_sb
g65871_da
g65871_db
g65871_sb
g65872_da
g65872_db
g65872_sb
g65875_da
g65875_db
g65875_sb
g65876_da
g65876_db
g65876_sb
g65877_da
g65877_db
g65877_sb
g65878_da
g65878_db
g65878_sb
g65882_da
g65882_db
g65882_sb
g65884_da
g65884_db
g65884_sb
g65885_da
g65885_db
g65885_sb
g65886_da
g65886_db
g65886_sb
g65890_da
g65890_db
g65890_sb
g65891_da
g65891_db
g65891_sb
g65892_da
g65892_db
g65892_sb
g65893_da
g65893_db
g65893_sb
g65894_da
g65894_db
g65894_sb
g65895_da
g65895_db
g65895_sb
g65896_da
g65896_db
g65896_sb
g65898_da
g65898_db
g65898_sb
g65899_da
g65899_db
g65899_sb
g65901_da
g65901_db
g65901_sb
g65902_da
g65902_db
g65902_sb
g65903_da
g65903_db
g65903_sb
g65904_da
g65904_db
g65904_sb
g65905_da
g65905_db
g65905_sb
g65907_da
g65907_db
g65907_sb
g65909_da
g65909_db
g65909_sb
g65910_da
g65910_db
g65910_sb
g65911_da
g65911_db
g65911_sb
g65912_da
g65912_db
g65912_sb
g65913_da
g65913_db
g65913_sb
g65915_da
g65915_db
g65915_sb
g65917_da
g65917_db
g65917_sb
g65918_da
g65918_db
g65918_sb
g65919_da
g65919_db
g65919_sb
g65920_da
g65920_db
g65920_sb
g65922_da
g65922_db
g65922_sb
g65923_da
g65923_db
g65923_sb
g65924_da
g65924_db
g65924_sb
g65926_da
g65926_db
g65926_sb
g65927_da
g65927_db
g65927_sb
g65929_da
g65929_db
g65930_da
g65930_db
g65930_sb
g65932_p
g65933_da
g65933_db
g65933_sb
g65934_da
g65934_db
g65934_sb
g65936_da
g65936_db
g65936_sb
g65937_p
g65938_p
g65939_p
g65940_da
g65940_db
g65940_sb
g65941_da
g65941_db
g65941_sb
g65942_da
g65942_db
g65942_sb
g65943_da
g65943_db
g65943_sb
g65944_da
g65944_db
g65944_sb
g65946_da
g65946_db
g65946_sb
g65947_da
g65947_db
g65947_sb
g65950_da
g65950_db
g65950_sb
g65951_da
g65951_db
g65951_sb
g65952_da
g65952_db
g65952_sb
g65954_da
g65954_db
g65954_sb
g65955_da
g65955_db
g65955_sb
g65956_da
g65956_db
g65956_sb
g65957_da
g65957_db
g65957_sb
g65958_da
g65958_db
g65958_sb
g65959_da
g65959_db
g65959_sb
g65960_da
g65960_db
g65960_sb
g65961_da
g65961_db
g65961_sb
g65962_da
g65962_db
g65962_sb
g65963_da
g65963_db
g65963_sb
g65967_da
g65967_db
g65967_sb
g65968_da
g65968_db
g65968_sb
g65969_da
g65969_db
g65969_sb
g65970_da
g65970_db
g65970_sb
g65971_da
g65971_db
g65971_sb
g65974_da
g65974_db
g65974_sb
g65975_da
g65975_db
g65975_sb
g65976_da
g65976_db
g65976_sb
g65977_da
g65977_db
g65977_sb
g65978_da
g65978_db
g65978_sb
g65982_p
g65983_p
g65984_p
g65985_p
g65986_p
g65988_p
g65989_p
g65990_p
g65992_p
g65993_p
g65994_da
g65994_db
g65994_sb
g65995_da
g65995_sb
g65996_da
g65996_sb
g65997_da
g65997_db
g65997_sb
g65998_da
g65998_db
g65999_da
g65999_db
g66001_sb
g66002_p
g66003_p
g66005_p
g66006_p
g66007_p
g66009_p
g66011_p
g66012_p
g66013_p
g66015_p
g66016_p
g66066_p
g66068_p
g66072_p
g66074_p
g66075_p
g66076_p
g66077_p
g66078_p
g66079_p
g66080_p
g66081_p
g66082_p
g66083_p
g66084_p
g66085_p
g66086_p
g66087_p
g66089_p
g66090_p
g66093_p
g66094_p
g66095_p
g66096_p
g66097_p
g66098_p
g66099_p
g66100_p
g66107_p
g66108_p
g66110_p
g66113_p
g66118_p
g66121_p
g66122_p
g66124_p
g66125_p
g66127_p
g66128_p
g66129_p
g66130_p
g66132_p
g66133_p
g66134_p
g66136_p
g66143_p
g66145_p
g66147_p
g66153_p
g66155_p
g66160_p
g66165_p
g66176_p
g66178_p
g66184_p
g66190_p
g66194_p
g66195_p
g66197_p
g66202_p
g66215_p
g66232_p
g66234_p
g66237_p
g66239_p
g66248_p
g66263_p
g66267_p
g66269_p
g66278_p
g66286_p
g66287_p
g66291_p
g66298_p
g66299_p
g66302_p
g66303_p
g66310_p
g66315_p
g66322_p
g66323_p
g66327_p
g66336_p
g66338_p
g66357_p
g66358_p
g66398_da
g66398_db
g66398_sb
g66399_da
g66399_db
g66399_sb
g66400_da
g66400_db
g66400_sb
g66401_da
g66401_db
g66401_sb
g66402_da
g66402_db
g66402_sb
g66403_da
g66403_db
g66403_sb
g66404_da
g66404_db
g66404_sb
g66406_da
g66406_db
g66407_da
g66407_db
g66407_sb
g66408_da
g66408_db
g66408_sb
g66409_da
g66409_db
g66409_sb
g66410_da
g66410_db
g66410_sb
g66411_da
g66411_db
g66411_sb
g66412_da
g66412_db
g66412_sb
g66413_da
g66413_db
g66413_sb
g66414_da
g66414_db
g66414_sb
g66415_da
g66415_db
g66415_sb
g66416_da
g66416_db
g66416_sb
g66417_da
g66417_db
g66417_sb
g66418_da
g66418_db
g66418_sb
g66419_da
g66419_db
g66419_sb
g66420_da
g66420_db
g66420_sb
g66421_da
g66421_db
g66422_da
g66422_db
g66422_sb
g66423_da
g66423_db
g66423_sb
g66424_da
g66424_db
g66424_sb
g66425_da
g66425_db
g66425_sb
g66426_da
g66426_db
g66426_sb
g66427_da
g66427_db
g66427_sb
g66428_da
g66428_db
g66428_sb
g66429_da
g66429_db
g66429_sb
g66430_da
g66430_db
g66430_sb
g66431_p
g66432_p
g66433_da
g66433_db
g66433_sb
g66434_p
g66435_p
g66436_p
g66437_p
g66438_p
g66439_p
g66443_p
g66444_p
g66447_p
g66450_p
g66452_p
g66453_p
g66455_p
g66456_da
g66456_db
g66456_sb
g66457_da
g66457_db
g66457_sb
g66458_p
g66458_p0
g66459_p
g66459_p0
g66464_p
g66464_p0
g66465_p
g66465_p0
g66473_p
g66475_p
g66477_da
g66477_db
g66477_sb
g66544_p
g66547_p
g66550_p
g66577_p
g66583_p
g66584_p
g66607_p
g66620_p
g66628_p
g66646_p
g66649_p
g66650_p
g66652_p
g66662_p
g66663_p
g66669_p
g66672_p
g66714_p
g66726_p
g66737_p
g66738_p
g66742_p
g66752_p
g66759_p
g66773_p
g66777_p
g66789_p
g66805_p
g66827_p
g66856_p
g66866_p
g66875_p
g66876_p
g66888_p
g66889_p
g66902_p
g66911_p
g66912_p
g66913_p
g66915_p
g66917_p
g66918_p
g66921_p
g66922_p
g66923_p
g66924_p
g66925_p
g66927_p
g66929_p
g66930_p
g66931_p
g66932_p
g66933_p
g66935_p
g66936_p
g66940_p
g66941_p
g66942_p
g66944_p
g66946_p
g66948_p
g66949_p
g66952_p
g66954_p
g66955_p
g66957_p
g66960_p
g66963_p
g66964_p
g66965_p
g66966_p
g66968_p
g66978_p
g66984_p
g66985_p
g66986_p
g66987_p
g66988_p
g66989_p
g66990_p
g66997_p
g67001_p
g67005_p
g67006_p
g67008_p
g67010_p
g67011_p
g67014_p
g67015_p
g67017_p
g67018_p
g67019_p
g67020_p
g67022_p
g67023_p
g67024_p
g67025_p
g67026_p
g67029_p
g67030_p
g67031_p
g67033_p
g67036_p
g67040_da
g67040_db
g67040_sb
g67041_da
g67041_db
g67042_da
g67042_db
g67042_sb
g67043_da
g67043_db
g67043_sb
g67044_da
g67044_db
g67044_sb
g67045_da
g67045_db
g67045_sb
g67046_da
g67046_db
g67046_sb
g67049_da
g67049_db
g67050_da
g67050_db
g67051_da
g67051_db
g67051_sb
g67052_db
g67053_da
g67053_db
g67053_sb
g67055_da
g67055_db
g67055_sb
g67056_da
g67056_db
g67058_da
g67058_db
g67059_da
g67059_db
g67067_da
g67067_db
g67068_da
g67068_db
g67069_da
g67069_db
g67071_da
g67071_db
g67071_sb
g67072_da
g67072_db
g67072_sb
g67073_da
g67073_db
g67074_da
g67074_db
g67075_da
g67075_db
g67083_da
g67083_db
g67084_da
g67084_db
g67084_sb
g67085_da
g67085_db
g67086_da
g67086_db
g67087_da
g67087_db
g67088_da
g67088_db
g67091_da
g67091_db
g67092_da
g67093_da
g67093_db
g67094_db
g67096_p
g67097_p
g67098_p
g67099_p
g67101_p
g67103_p
g67104_p
g67105_p
g67106_p
g67107_p
g67108_p
g67109_p
g67110_p
g67111_p
g67112_p
g67113_p
g67114_p
g67115_p
g67116_p
g67117_p
g67118_p
g67119_p
g67120_p
g67122_p
g67123_p
g67124_p
g67125_p
g67126_p
g67127_p
g67128_p
g67129_p
g67130_p
g67131_p
g67133_p
g67134_p
g67135_p
g67137_p
g67138_p
g67139_p
g67140_p
g67141_p
g67143_p
g67144_p
g67147_p
g67148_p
g67149_p
g67150_p
g67151_p
g67152_p
g67153_p
g67154_p
g67155_p
g67157_p
g67311_p
g67324_p
g67327_p
g67340_p
g67353_p
g67355_p
g67364_p
g67371_p
g67386_p
g67389_p
g67392_p
g67396_p
g67397_p
g67405_p
g67411_p
g67421_p
g67425_p
g67430_p
g67432_p
g67434_p
g67437_p
g67446_p
g67453_p
g67457_p
g67459_p
g67468_p
g67498_p
g67502_p
g67506_p
g67507_p
g67523_p
g67531_p
g67534_p
g67535_p
g67537_p
g67538_p
g67544_p
g67549_p
g67559_p
g67581_p
g67582_p
g67583_p
g67592_p
g67600_p
g67603_p
g67610_p
g67624_p
g67625_p
g67626_p
g67631_p
g67671_p
g67672_p
g67675_p
g67680_p
g67688_p
g67689_p
g67699_p
g67712_p
g67721_p
g67725_p
g67731_p
g67735_p
g67739_p
g67740_p
g67746_p
g67747_p
g67754_p
g67757_p
g67758_p
g67763_p
g67778_p
g67791_p
g67799_p
g67802_p
g67804_p
g67806_p
g67807_p
g67814_p
g67828_p
g68_p
g73989_p
g74028_p
g74116_dup_p
g74118_p
g74140_p
g74153_p
g74162_dup_p
g74174_p
g74243_p
g74245_p
g74270_p
g74283_p
g74363_p
g74408_p
g74429_p
g74509_p
g74510_p
g74553_p
g74563_p
g74567_p
g74576_p
g74580_p
g74630_p
g74644_p
g74671_p
g74689_p
g74739_p
g74787_p
g74879_p
g74920_p
g74930_p
g74956_p
g74958_p1
g74958_p2
g74981_p
g74982_p
g74998_da
g74998_db
g74998_sb
g75024_da
g75024_db
g75024_sb
g75059_p
g75072_da
g75088_p
g75091_da
g75091_db
g75091_sb
g75126_p
g75129_p
g75160_da
g75160_db
g75160_sb
g75162_da
g75162_db
g75162_sb
g75177_da
g75177_db
g75177_sb
g75178_da
g75178_db
g75178_sb
g75181_da
g75181_db
g75181_sb
g75202_da
g75202_db
g75202_sb
g75413_da
g75413_db
g75413_sb
g75416_da
g75416_db
g75416_sb
g75418_da
g75418_db
g75418_sb
g75_p
i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_29__Q
i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_31__Q
i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_0__Q
i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_10__Q
i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_11__Q
i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_12__Q
i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_13__Q
i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_14__Q
i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_15__Q
i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_16__Q
i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_17__Q
i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_18__Q
i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_19__Q
i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_1__Q
i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_20__Q
i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_21__Q
i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_22__Q
i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_23__Q
i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_24__Q
i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_25__Q
i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_26__Q
i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_27__Q
i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_28__Q
i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_29__Q
i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_2__Q
i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_30__Q
i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_31__Q
i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_3__Q
i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_4__Q
i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_5__Q
i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_6__Q
i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_7__Q
i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_8__Q
i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_9__Q
i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid
n_10002
n_1001
n_10010
n_10014
n_10017
n_10020
n_10023
n_10026
n_10029
n_10032
n_10035
n_10038
n_10048
n_1005
n_10051
n_10054
n_10057
n_10060
n_10063
n_10066
n_10069
n_1007
n_10078
n_1008
n_10087
n_1009
n_10090
n_10093
n_10096
n_10099
n_10102
n_10105
n_10106
n_10112
n_10113
n_10116
n_10117
n_1012
n_10120
n_10121
n_10124
n_10127
n_10128
n_1013
n_10131
n_10134
n_10135
n_10139
n_1014
n_10141
n_10144
n_10147
n_10148
n_10151
n_10154
n_10157
n_1016
n_10160
n_10163
n_10168
n_1017
n_10170
n_10173
n_10176
n_10179
n_10180
n_10183
n_10185
n_10188
n_1019
n_10190
n_10195
n_10198
n_10199
n_10202
n_10205
n_10206
n_10213
n_10216
n_1022
n_10221
n_10225
n_1023
n_10232
n_10235
n_10236
n_10237
n_1024
n_10244
n_10247
n_1025
n_10250
n_10256
n_10257
n_10258
n_1026
n_10261
n_10263
n_1027
n_10270
n_10272
n_10274
n_10275
n_10276
n_10277
n_10278
n_10279
n_1028
n_10281
n_10286
n_10288
n_1029
n_10291
n_10294
n_10304
n_10306
n_1031
n_10310
n_10314
n_10316
n_10317
n_10319
n_1032
n_10321
n_10323
n_10325
n_10327
n_10329
n_1033
n_10331
n_10332
n_10334
n_10336
n_10338
n_1034
n_10340
n_10342
n_10344
n_10348
n_10349
n_1035
n_10351
n_10353
n_1036
n_10361
n_10362
n_10363
n_10365
n_10366
n_1037
n_10370
n_10376
n_10377
n_10378
n_1038
n_10380
n_10381
n_10383
n_10385
n_1039
n_10390
n_10393
n_10394
n_10397
n_10399
n_10400
n_10401
n_10402
n_10404
n_10405
n_10408
n_1041
n_10410
n_10411
n_10412
n_10413
n_10414
n_10416
n_10418
n_10419
n_10421
n_10423
n_10424
n_10426
n_10428
n_10432
n_10436
n_10438
n_10440
n_10441
n_10444
n_10446
n_10449
n_10450
n_10453
n_10455
n_10457
n_10459
n_10460
n_10462
n_10464
n_10465
n_10467
n_10469
n_10470
n_10474
n_10476
n_10477
n_10478
n_10479
n_10481
n_10483
n_10485
n_10487
n_10489
n_10491
n_10493
n_10495
n_10497
n_10501
n_10506
n_10508
n_10511
n_10513
n_10518
n_10521
n_10524
n_10527
n_10530
n_10538
n_10541
n_10544
n_10553
n_10554
n_10556
n_10559
n_10560
n_10566
n_10569
n_1057
n_10572
n_10575
n_10584
n_10588
n_10592
n_10595
n_10596
n_10599
n_10602
n_10605
n_10608
n_1061
n_10611
n_10614
n_10617
n_10624
n_10627
n_1063
n_10630
n_10634
n_10637
n_10638
n_1064
n_10641
n_10644
n_10647
n_10650
n_10653
n_10656
n_10659
n_10660
n_10661
n_10662
n_10669
n_10672
n_10675
n_10676
n_10679
n_10680
n_10681
n_10685
n_10688
n_1069
n_10691
n_10693
n_10696
n_10708
n_10711
n_10715
n_1072
n_10728
n_1073
n_10731
n_10734
n_10738
n_1074
n_10741
n_10744
n_10747
n_10750
n_10753
n_10754
n_10755
n_10758
n_10763
n_10764
n_10765
n_10768
n_1077
n_10771
n_10774
n_10784
n_10785
n_10787
n_10788
n_10789
n_1079
n_10791
n_10792
n_10793
n_10795
n_10799
n_1080
n_10802
n_10803
n_10804
n_10807
n_1081
n_10813
n_10815
n_10820
n_10821
n_10825
n_10828
n_10829
n_1083
n_10832
n_10833
n_10834
n_10835
n_10836
n_10839
n_10843
n_10847
n_10848
n_1085
n_10851
n_10853
n_10856
n_10859
n_1086
n_10860
n_10865
n_10866
n_10867
n_10870
n_10873
n_10875
n_10876
n_10877
n_10881
n_10885
n_1089
n_10892
n_10901
n_10902
n_10904
n_10905
n_10906
n_10909
n_1091
n_10912
n_10913
n_10916
n_10917
n_10919
n_10922
n_10923
n_10927
n_1093
n_10930
n_10931
n_10932
n_10936
n_10939
n_1094
n_10942
n_10944
n_1095
n_10951
n_10952
n_10956
n_1096
n_10961
n_10962
n_10963
n_10967
n_10970
n_10971
n_10974
n_10975
n_10976
n_10977
n_10978
n_10981
n_10985
n_10986
n_10987
n_1099
n_10991
n_11
n_1100
n_11002
n_11005
n_11008
n_1101
n_11013
n_11014
n_11019
n_1103
n_11034
n_11036
n_11037
n_11038
n_1104
n_11040
n_11041
n_11044
n_11046
n_11047
n_11048
n_11049
n_11050
n_11051
n_11053
n_11054
n_11055
n_11056
n_11057
n_11058
n_11059
n_11060
n_11061
n_11062
n_11065
n_11066
n_11069
n_1107
n_11070
n_11071
n_11072
n_11073
n_1108
n_11083
n_11084
n_11085
n_11086
n_11087
n_11088
n_11089
n_1109
n_11090
n_11094
n_11095
n_11096
n_11097
n_11099
n_1110
n_11100
n_11101
n_11102
n_11104
n_11106
n_11107
n_11108
n_11109
n_1111
n_11110
n_11111
n_11113
n_11115
n_11118
n_11119
n_11120
n_11121
n_11122
n_11123
n_11124
n_11125
n_11126
n_11129
n_11130
n_11131
n_11132
n_11134
n_11135
n_11136
n_11137
n_11138
n_11139
n_11140
n_11142
n_11143
n_11144
n_11145
n_11146
n_11148
n_11149
n_1115
n_11152
n_11157
n_11158
n_1116
n_11162
n_11164
n_11165
n_11169
n_1117
n_11174
n_11175
n_11177
n_11178
n_11179
n_1118
n_11180
n_11181
n_11182
n_11184
n_11188
n_1119
n_11190
n_11191
n_11198
n_112
n_11202
n_11203
n_11205
n_11206
n_11207
n_11208
n_11211
n_11212
n_11213
n_11214
n_11215
n_11216
n_11217
n_11218
n_11219
n_1122
n_11220
n_11223
n_11224
n_11226
n_11228
n_1123
n_11232
n_11234
n_11236
n_11238
n_11239
n_1124
n_11240
n_11242
n_11243
n_11244
n_11245
n_11246
n_11247
n_11249
n_1125
n_11250
n_11251
n_11252
n_11254
n_11255
n_11259
n_11261
n_11264
n_11265
n_11266
n_11268
n_11270
n_11271
n_11273
n_11274
n_11276
n_11277
n_11279
n_11280
n_11281
n_11282
n_11283
n_11284
n_11285
n_11289
n_11290
n_11293
n_11295
n_11297
n_11302
n_11305
n_11306
n_11307
n_11309
n_11311
n_11314
n_11318
n_11320
n_11322
n_11324
n_11326
n_11327
n_11328
n_1133
n_11330
n_11332
n_11334
n_11337
n_11338
n_1134
n_11340
n_11342
n_11344
n_11345
n_11347
n_11349
n_1135
n_11350
n_11352
n_11353
n_11355
n_11357
n_1136
n_11361
n_11362
n_11363
n_11365
n_11367
n_11369
n_1137
n_11370
n_11372
n_11373
n_11375
n_11377
n_11379
n_1138
n_11380
n_11383
n_11385
n_11386
n_11388
n_1139
n_11390
n_11391
n_11393
n_11396
n_11398
n_11399
n_11403
n_11405
n_11406
n_11408
n_11410
n_11411
n_11414
n_11415
n_11417
n_11418
n_11419
n_1142
n_11420
n_11421
n_11423
n_11424
n_11425
n_11427
n_11429
n_1143
n_11432
n_11434
n_11435
n_11436
n_11437
n_11438
n_11440
n_11441
n_11445
n_11446
n_11448
n_11449
n_1145
n_11450
n_11452
n_11456
n_11457
n_11458
n_1146
n_11460
n_11462
n_11463
n_11464
n_11467
n_1147
n_11470
n_11472
n_11473
n_11474
n_11476
n_11477
n_11479
n_11480
n_11483
n_11484
n_11487
n_11489
n_11490
n_11492
n_11495
n_11496
n_11497
n_11499
n_1150
n_11500
n_11505
n_11507
n_11509
n_1151
n_11512
n_11513
n_11515
n_11516
n_11517
n_11519
n_1152
n_11521
n_11523
n_11524
n_11526
n_11528
n_1153
n_11530
n_11531
n_11532
n_11533
n_11535
n_11536
n_1154
n_11540
n_11542
n_11543
n_11544
n_11545
n_11546
n_11547
n_11548
n_1155
n_11553
n_11556
n_11557
n_11559
n_11560
n_11562
n_11564
n_11565
n_11566
n_11568
n_1157
n_11570
n_11572
n_11573
n_11579
n_11582
n_11584
n_11585
n_11586
n_11587
n_11588
n_11589
n_1159
n_11590
n_11593
n_11595
n_11597
n_11598
n_1160
n_11601
n_11603
n_11605
n_11606
n_11609
n_1161
n_11613
n_11614
n_11616
n_11617
n_11618
n_1162
n_11620
n_11622
n_11623
n_11624
n_11625
n_11626
n_11630
n_11633
n_11634
n_11635
n_11637
n_11638
n_1164
n_11640
n_11642
n_11644
n_11648
n_1165
n_11650
n_11651
n_11652
n_11653
n_11655
n_11657
n_11659
n_1166
n_11660
n_11661
n_11663
n_11665
n_11666
n_11667
n_11668
n_11669
n_1167
n_11670
n_11671
n_11674
n_11679
n_1168
n_11680
n_11681
n_11682
n_11683
n_11685
n_11686
n_11687
n_11688
n_11689
n_1169
n_11690
n_11692
n_11694
n_11695
n_11697
n_11698
n_1170
n_11701
n_11703
n_11708
n_11710
n_11716
n_11717
n_11719
n_11723
n_11725
n_11728
n_1173
n_11730
n_11732
n_11734
n_11735
n_11736
n_11739
n_1174
n_11740
n_11741
n_11744
n_1176
n_11762
n_11767
n_1177
n_11773
n_11775
n_11776
n_11777
n_11781
n_11782
n_11783
n_11784
n_11786
n_11788
n_11790
n_11791
n_11792
n_11793
n_11795
n_11799
n_1180
n_11803
n_11804
n_11807
n_11808
n_11809
n_11810
n_11811
n_11815
n_11816
n_11817
n_11818
n_11820
n_11821
n_11822
n_11824
n_11825
n_11826
n_11827
n_11829
n_1183
n_11830
n_11831
n_11832
n_11833
n_11834
n_11835
n_11836
n_11840
n_11844
n_11845
n_11846
n_11847
n_11848
n_11849
n_1185
n_11850
n_11851
n_11852
n_11853
n_11854
n_11855
n_11856
n_11857
n_11858
n_11859
n_1186
n_11860
n_11861
n_11862
n_11863
n_11864
n_11865
n_11866
n_11867
n_11868
n_11869
n_1187
n_11870
n_11871
n_11872
n_11873
n_11874
n_11875
n_11876
n_11877
n_11878
n_1188
n_11880
n_11881
n_11884
n_11886
n_11887
n_1189
n_11890
n_11893
n_11897
n_11898
n_11899
n_119
n_1190
n_11900
n_11901
n_11902
n_11907
n_11910
n_11911
n_11917
n_11920
n_11921
n_11922
n_11923
n_11927
n_11928
n_11929
n_11930
n_11934
n_11935
n_11936
n_11940
n_11945
n_11950
n_11951
n_11952
n_1196
n_11968
n_1197
n_11970
n_11975
n_11977
n_11979
n_1198
n_11982
n_11986
n_11987
n_11988
n_1199
n_11991
n_11999
n_12
n_1200
n_12000
n_12001
n_12002
n_12004
n_12007
n_12008
n_1201
n_12010
n_12011
n_12012
n_12013
n_12019
n_12020
n_12021
n_12022
n_12023
n_12026
n_12030
n_12035
n_12036
n_12037
n_12038
n_1204
n_12040
n_12041
n_12042
n_12046
n_12049
n_12050
n_12052
n_12053
n_12054
n_12055
n_12056
n_12057
n_12060
n_12062
n_12064
n_12065
n_12066
n_12069
n_1207
n_12071
n_12078
n_1208
n_12081
n_12084
n_12085
n_12087
n_12088
n_12089
n_1209
n_12090
n_12091
n_12092
n_12095
n_12097
n_12098
n_12099
n_12100
n_12101
n_12102
n_12103
n_12105
n_12109
n_1211
n_12114
n_12115
n_12116
n_12118
n_12121
n_12124
n_12125
n_12128
n_12129
n_1213
n_12132
n_12133
n_12134
n_12135
n_12137
n_12139
n_12140
n_12141
n_12143
n_12144
n_12145
n_12147
n_12148
n_1215
n_12151
n_12153
n_12154
n_12155
n_12156
n_12158
n_12159
n_1216
n_12160
n_12161
n_12162
n_12163
n_12164
n_12165
n_12166
n_12167
n_12168
n_12169
n_1217
n_12170
n_12179
n_1218
n_12181
n_12183
n_12184
n_12185
n_12186
n_12187
n_12188
n_1219
n_12190
n_12191
n_12192
n_12196
n_12198
n_12199
n_1220
n_12200
n_1221
n_12210
n_12211
n_12214
n_12215
n_12216
n_12217
n_12218
n_12220
n_12221
n_12222
n_12223
n_12225
n_12226
n_12227
n_12228
n_12229
n_12230
n_12232
n_12233
n_12234
n_12237
n_12238
n_12239
n_1224
n_12241
n_12242
n_12243
n_12244
n_1225
n_12251
n_12255
n_12256
n_12257
n_12258
n_12264
n_12265
n_12266
n_12267
n_12268
n_12269
n_1227
n_12270
n_12271
n_12272
n_12273
n_12274
n_12276
n_12277
n_1228
n_12280
n_12282
n_12283
n_12287
n_12289
n_1229
n_12290
n_12291
n_12292
n_12293
n_12294
n_12297
n_123
n_12300
n_12301
n_12307
n_12309
n_1231
n_12310
n_12312
n_12313
n_12314
n_12319
n_12320
n_12322
n_12327
n_12328
n_12329
n_12330
n_12333
n_12334
n_12344
n_12346
n_12350
n_12351
n_12354
n_12355
n_12356
n_12357
n_12358
n_12359
n_12362
n_12363
n_12364
n_12367
n_12369
n_12370
n_12371
n_12372
n_12373
n_12374
n_12377
n_1238
n_12381
n_12382
n_12383
n_12385
n_12386
n_12388
n_12389
n_12390
n_12391
n_12394
n_12396
n_12398
n_12401
n_12403
n_12404
n_12405
n_12406
n_12408
n_1241
n_12410
n_12411
n_12412
n_12413
n_12417
n_1242
n_12420
n_12422
n_12423
n_12424
n_12425
n_12426
n_12427
n_12429
n_12430
n_12432
n_12433
n_12434
n_12438
n_12439
n_12440
n_12441
n_12449
n_12451
n_12453
n_12455
n_12458
n_12459
n_12461
n_12462
n_12464
n_12465
n_12466
n_12468
n_12469
n_12470
n_12471
n_12472
n_12473
n_12474
n_12476
n_12478
n_1248
n_12483
n_12485
n_12486
n_12487
n_12491
n_12492
n_12493
n_12494
n_12502
n_12506
n_12509
n_1251
n_12510
n_12511
n_12512
n_12513
n_12514
n_12515
n_12516
n_12518
n_1252
n_12520
n_12522
n_12523
n_12524
n_12526
n_12527
n_12529
n_1253
n_12530
n_12531
n_12532
n_12533
n_12534
n_12535
n_12536
n_12537
n_12538
n_12539
n_12540
n_12541
n_12542
n_12543
n_12544
n_12545
n_12546
n_12547
n_12548
n_12549
n_12550
n_12551
n_12552
n_12553
n_12554
n_12555
n_12556
n_12557
n_12558
n_12559
n_12560
n_12561
n_12562
n_12563
n_12565
n_12566
n_12568
n_12569
n_12570
n_12571
n_12572
n_12573
n_12574
n_12575
n_12577
n_12578
n_12579
n_1258
n_12580
n_12581
n_12583
n_12584
n_12585
n_12586
n_12587
n_12588
n_12589
n_1259
n_12590
n_12591
n_12595
n_12599
n_1260
n_12600
n_12602
n_12603
n_12606
n_12607
n_1261
n_12612
n_12617
n_12619
n_12620
n_12621
n_12622
n_12628
n_12629
n_1263
n_12630
n_12631
n_12632
n_12633
n_12634
n_12638
n_12639
n_1264
n_12640
n_12641
n_12642
n_12643
n_12645
n_12646
n_12647
n_12648
n_12649
n_1265
n_12650
n_12651
n_12653
n_12655
n_12656
n_12658
n_12659
n_1266
n_12661
n_12662
n_12665
n_12668
n_12669
n_12670
n_12671
n_12672
n_12673
n_12674
n_12680
n_12685
n_12686
n_12687
n_1269
n_12690
n_12693
n_12695
n_12696
n_12697
n_12699
n_1270
n_12700
n_12701
n_12702
n_12703
n_12704
n_12705
n_12706
n_12707
n_12709
n_1271
n_12710
n_12711
n_12714
n_12715
n_12716
n_12717
n_1272
n_12721
n_12722
n_12723
n_12725
n_12726
n_12727
n_12728
n_12729
n_1273
n_12731
n_12732
n_12734
n_12736
n_12737
n_12738
n_1274
n_12741
n_12744
n_12745
n_12746
n_12747
n_12748
n_12749
n_1275
n_12754
n_12756
n_1276
n_12760
n_12761
n_12762
n_12763
n_12765
n_12768
n_12769
n_1277
n_12770
n_12771
n_12772
n_12773
n_12774
n_12775
n_12781
n_12784
n_12786
n_12787
n_12788
n_12789
n_1279
n_12791
n_12797
n_12798
n_12799
n_1280
n_12801
n_12805
n_12806
n_1281
n_12811
n_12813
n_12815
n_12816
n_12817
n_12818
n_12819
n_1282
n_12821
n_12822
n_12823
n_12824
n_12825
n_12826
n_12827
n_1283
n_12830
n_12831
n_12833
n_12834
n_12835
n_12836
n_12837
n_12839
n_1284
n_12840
n_12841
n_12842
n_12843
n_12845
n_12846
n_12847
n_12848
n_12849
n_1285
n_12850
n_12851
n_12852
n_12853
n_12855
n_12858
n_1286
n_12862
n_12864
n_12865
n_12866
n_12870
n_12871
n_12872
n_12873
n_12878
n_12879
n_1288
n_12880
n_12881
n_12883
n_12884
n_12885
n_12886
n_12887
n_12888
n_12889
n_1289
n_12890
n_12892
n_12893
n_12894
n_12896
n_12897
n_12898
n_12899
n_1290
n_12900
n_12901
n_12902
n_12903
n_12907
n_1291
n_12914
n_12915
n_12916
n_12917
n_12918
n_12919
n_12920
n_12921
n_12922
n_12924
n_12928
n_12929
n_1293
n_12930
n_12931
n_12932
n_12933
n_12934
n_12936
n_12937
n_1294
n_12940
n_12941
n_12942
n_12947
n_12948
n_12951
n_12952
n_12954
n_12956
n_12957
n_12958
n_12959
n_12961
n_12962
n_12963
n_12966
n_12968
n_12970
n_12972
n_12974
n_12976
n_12978
n_12980
n_12981
n_12982
n_12983
n_12984
n_12985
n_12986
n_12988
n_1299
n_12990
n_12992
n_12994
n_12996
n_12998
n_13000
n_13002
n_13004
n_13006
n_13008
n_13010
n_13012
n_13014
n_13016
n_13018
n_13020
n_13022
n_13024
n_13026
n_13027
n_13028
n_13036
n_1304
n_13041
n_13043
n_13045
n_13046
n_13047
n_13050
n_13052
n_13054
n_13056
n_13058
n_13059
n_1306
n_13060
n_13061
n_13065
n_13066
n_13073
n_13074
n_13075
n_13076
n_13077
n_13078
n_13079
n_13080
n_13081
n_13082
n_13083
n_13084
n_13085
n_13086
n_13087
n_13088
n_13089
n_13090
n_13091
n_13093
n_13094
n_13095
n_13097
n_13098
n_13100
n_13102
n_13104
n_13105
n_13106
n_13107
n_13111
n_13113
n_13115
n_13116
n_13120
n_13122
n_13123
n_13124
n_13125
n_13127
n_13128
n_13129
n_13130
n_13131
n_13132
n_13133
n_13134
n_13135
n_13137
n_13138
n_13139
n_13140
n_13141
n_13142
n_13143
n_13144
n_13145
n_13148
n_1315
n_13150
n_13152
n_13155
n_13157
n_1316
n_13160
n_13164
n_13165
n_13167
n_13169
n_1317
n_13170
n_13171
n_13173
n_13175
n_13176
n_13178
n_13179
n_1318
n_13180
n_13181
n_13182
n_13184
n_13185
n_13186
n_13187
n_13189
n_13190
n_13191
n_13192
n_13195
n_13197
n_13199
n_13200
n_13201
n_13203
n_13205
n_13208
n_13210
n_13211
n_13213
n_13214
n_13215
n_13217
n_1322
n_13220
n_13221
n_13222
n_13223
n_13228
n_13231
n_13235
n_13239
n_13241
n_13244
n_13246
n_13249
n_1325
n_13251
n_13254
n_13256
n_13258
n_1326
n_13260
n_13263
n_13266
n_13271
n_13273
n_13275
n_13277
n_13279
n_13281
n_13283
n_13284
n_13285
n_13286
n_13287
n_1329
n_13292
n_13294
n_13295
n_1330
n_13302
n_13303
n_13304
n_13305
n_13306
n_13308
n_1331
n_13311
n_13313
n_13315
n_13318
n_1332
n_13320
n_13321
n_13323
n_13326
n_13328
n_1333
n_13331
n_13334
n_13336
n_13337
n_13338
n_13339
n_1334
n_13340
n_13341
n_13342
n_13343
n_13344
n_13345
n_13348
n_13349
n_1335
n_13350
n_13351
n_13353
n_13354
n_13355
n_13356
n_13357
n_13358
n_13359
n_1336
n_13360
n_13361
n_13362
n_13363
n_13365
n_13366
n_13368
n_13369
n_1337
n_13370
n_13371
n_13372
n_13373
n_13374
n_13375
n_13376
n_13378
n_13379
n_1338
n_13380
n_13381
n_13383
n_13384
n_13386
n_13387
n_13388
n_13389
n_13390
n_13391
n_13392
n_13393
n_13394
n_13395
n_13398
n_13399
n_1340
n_13400
n_13401
n_13402
n_13403
n_13404
n_13405
n_13406
n_13407
n_13408
n_13409
n_1341
n_13410
n_13411
n_13412
n_13413
n_13414
n_13415
n_13416
n_13417
n_13418
n_13419
n_1342
n_13420
n_13421
n_13422
n_13423
n_13424
n_13425
n_13426
n_13427
n_13428
n_13429
n_1343
n_13430
n_13431
n_13432
n_13434
n_13435
n_13436
n_13437
n_13438
n_13439
n_1344
n_13441
n_13442
n_13444
n_13445
n_13446
n_13447
n_13448
n_13449
n_1345
n_13450
n_13452
n_13453
n_13454
n_13455
n_13457
n_13459
n_1346
n_13461
n_13462
n_13463
n_13464
n_13466
n_13467
n_13468
n_13469
n_1347
n_13470
n_13474
n_13475
n_13481
n_13482
n_13483
n_13484
n_13485
n_13486
n_13487
n_13488
n_13489
n_1349
n_13490
n_13493
n_13495
n_13496
n_13497
n_135
n_1350
n_13500
n_13503
n_13504
n_13505
n_13506
n_13508
n_13509
n_1351
n_13511
n_13512
n_13516
n_13517
n_13518
n_13519
n_1352
n_13520
n_13522
n_13523
n_13524
n_13526
n_13528
n_13529
n_1353
n_13531
n_13532
n_13533
n_13534
n_13535
n_13536
n_13538
n_13539
n_1354
n_13540
n_13544
n_13546
n_13547
n_1355
n_13552
n_13556
n_13557
n_13558
n_13559
n_1356
n_13560
n_13561
n_13562
n_13563
n_13565
n_13566
n_13567
n_13568
n_1357
n_13570
n_13573
n_13574
n_13575
n_13576
n_13577
n_1358
n_13581
n_13582
n_13583
n_13584
n_13585
n_13587
n_13589
n_1359
n_13591
n_13592
n_13593
n_13595
n_13597
n_13599
n_1360
n_13601
n_13603
n_13605
n_13607
n_13608
n_13609
n_1361
n_13610
n_13611
n_13613
n_13614
n_13616
n_13617
n_13618
n_13619
n_1362
n_13620
n_13621
n_13622
n_13623
n_13624
n_13625
n_13628
n_13629
n_1363
n_13631
n_13632
n_13634
n_13635
n_13636
n_13638
n_1364
n_13640
n_13641
n_13642
n_13643
n_13645
n_13646
n_13647
n_13648
n_13649
n_1365
n_13650
n_13651
n_13652
n_13653
n_13654
n_13655
n_13657
n_13658
n_13659
n_1366
n_13661
n_13662
n_13663
n_13664
n_13665
n_13666
n_13668
n_13669
n_13670
n_13671
n_13672
n_13673
n_13674
n_13678
n_13679
n_13680
n_13681
n_13682
n_13685
n_13686
n_13687
n_13688
n_1369
n_13691
n_13694
n_13695
n_13696
n_13697
n_13698
n_1370
n_13701
n_13704
n_13705
n_13709
n_1371
n_13710
n_13711
n_13712
n_13717
n_13719
n_1372
n_13720
n_13721
n_13722
n_13724
n_13725
n_13727
n_13728
n_13729
n_13731
n_13732
n_13734
n_13735
n_13736
n_13738
n_13740
n_13741
n_13743
n_13744
n_13745
n_13747
n_13748
n_13749
n_1375
n_13754
n_13755
n_13756
n_13757
n_13759
n_1376
n_13760
n_13761
n_13762
n_13763
n_13764
n_13766
n_1377
n_13770
n_13771
n_13772
n_13773
n_13776
n_13777
n_13778
n_1378
n_13780
n_13783
n_13784
n_13785
n_13786
n_13787
n_13789
n_1379
n_13790
n_13792
n_13793
n_13794
n_13798
n_1380
n_13800
n_13806
n_13807
n_13809
n_1381
n_13810
n_13812
n_13813
n_13814
n_13815
n_13816
n_13817
n_13819
n_1382
n_13820
n_13821
n_13822
n_13823
n_13825
n_13827
n_13828
n_13829
n_1383
n_13830
n_1384
n_13842
n_13843
n_13844
n_13845
n_13847
n_1385
n_13850
n_13851
n_13854
n_13856
n_13857
n_13859
n_13862
n_13864
n_13866
n_13867
n_13869
n_1387
n_13870
n_13871
n_13872
n_13873
n_13874
n_13875
n_13876
n_13878
n_1388
n_13880
n_13881
n_13882
n_13885
n_13886
n_13888
n_13889
n_1389
n_13891
n_13895
n_13896
n_13898
n_139
n_1390
n_13901
n_13905
n_13907
n_13908
n_1391
n_13910
n_13911
n_13917
n_13919
n_1392
n_13920
n_13921
n_13922
n_13924
n_1393
n_13935
n_13936
n_13937
n_13938
n_13939
n_1394
n_13940
n_13941
n_13942
n_13943
n_13944
n_13945
n_13948
n_1395
n_13951
n_13952
n_13953
n_13954
n_13955
n_13957
n_13959
n_1396
n_13960
n_13961
n_13966
n_13967
n_13968
n_1397
n_13971
n_13972
n_13973
n_13974
n_13976
n_13977
n_13980
n_13983
n_13984
n_13987
n_1399
n_13990
n_13991
n_13993
n_13995
n_13996
n_13998
n_14
n_14001
n_14008
n_14009
n_1401
n_14011
n_14012
n_14013
n_14014
n_14015
n_14017
n_14019
n_1402
n_14020
n_14021
n_14023
n_14024
n_14025
n_14026
n_14027
n_14029
n_14030
n_14031
n_14033
n_14035
n_14037
n_14038
n_14039
n_1404
n_14042
n_14043
n_14045
n_14046
n_14049
n_1405
n_14050
n_14056
n_14057
n_1406
n_14060
n_14068
n_14069
n_1407
n_14070
n_14072
n_14073
n_14074
n_14075
n_14076
n_14077
n_14078
n_14079
n_1408
n_14080
n_14081
n_14082
n_14083
n_14084
n_14085
n_14086
n_14087
n_14088
n_1409
n_14091
n_14092
n_14093
n_14094
n_14095
n_14096
n_14098
n_1410
n_14103
n_14104
n_14105
n_14106
n_14107
n_14108
n_14109
n_1411
n_14110
n_14111
n_14112
n_14113
n_14114
n_14115
n_14116
n_14117
n_14118
n_1412
n_14120
n_14125
n_14126
n_14127
n_14128
n_1413
n_14132
n_14133
n_14134
n_14138
n_1414
n_14140
n_1415
n_14154
n_14155
n_14160
n_14161
n_14163
n_14166
n_14167
n_14170
n_14171
n_14172
n_14175
n_14176
n_14177
n_14178
n_14179
n_1418
n_14180
n_14182
n_14184
n_14185
n_14186
n_14187
n_14188
n_14189
n_1419
n_14190
n_14191
n_14192
n_14193
n_14194
n_14195
n_14196
n_14197
n_14198
n_14199
n_1420
n_14200
n_14206
n_14207
n_1421
n_14213
n_14214
n_14216
n_14218
n_1422
n_14220
n_14222
n_14227
n_14228
n_14229
n_1423
n_14230
n_1424
n_14246
n_14247
n_1425
n_14251
n_14252
n_14253
n_14255
n_14256
n_1426
n_14261
n_14263
n_14264
n_14267
n_14268
n_14269
n_14270
n_14273
n_14274
n_14275
n_14276
n_1428
n_14283
n_14284
n_1429
n_14296
n_14297
n_143
n_14300
n_14303
n_14304
n_14305
n_14306
n_14307
n_14309
n_1431
n_14311
n_14313
n_14314
n_14315
n_14317
n_1432
n_14323
n_14324
n_14325
n_14326
n_14327
n_14328
n_14329
n_1433
n_14330
n_14331
n_14332
n_14333
n_14334
n_14335
n_14336
n_14337
n_14338
n_14339
n_1434
n_14340
n_14341
n_14342
n_14343
n_14344
n_14345
n_14346
n_14349
n_1435
n_14350
n_14351
n_14353
n_14354
n_14355
n_14356
n_14357
n_14358
n_14359
n_1436
n_14360
n_14361
n_14362
n_14363
n_14367
n_14368
n_14369
n_1437
n_14370
n_14371
n_14372
n_14375
n_14379
n_1438
n_14380
n_14381
n_14382
n_14383
n_14384
n_14385
n_14389
n_14399
n_1440
n_14402
n_14403
n_14407
n_14408
n_1441
n_14410
n_14413
n_14414
n_14415
n_14416
n_14419
n_1442
n_14420
n_14421
n_14422
n_14428
n_14429
n_1443
n_14430
n_14431
n_14432
n_14433
n_14434
n_14436
n_14437
n_14438
n_14439
n_1444
n_14440
n_14441
n_14442
n_14443
n_14448
n_14449
n_1445
n_14450
n_14451
n_14454
n_14455
n_14456
n_14457
n_14458
n_1446
n_14460
n_14461
n_14467
n_1447
n_14472
n_14478
n_14479
n_1448
n_14482
n_14483
n_14484
n_14485
n_14486
n_14487
n_14489
n_1449
n_14491
n_14494
n_14495
n_14497
n_14498
n_14500
n_14504
n_14505
n_14506
n_14507
n_14508
n_14511
n_14512
n_14513
n_14514
n_14515
n_14516
n_14517
n_14518
n_14519
n_1452
n_14521
n_14526
n_14527
n_14528
n_14529
n_1453
n_14530
n_14532
n_14534
n_14535
n_14536
n_14539
n_1454
n_14541
n_14544
n_14545
n_14546
n_14547
n_14548
n_14550
n_14554
n_14556
n_14557
n_14559
n_14560
n_14567
n_14570
n_14571
n_14576
n_14578
n_14579
n_14582
n_14583
n_14585
n_14588
n_14589
n_14590
n_14591
n_14593
n_14594
n_14595
n_14596
n_14598
n_14599
n_1460
n_14601
n_14602
n_14603
n_14604
n_14605
n_14607
n_14608
n_1461
n_14610
n_14611
n_14612
n_14613
n_14614
n_14615
n_14616
n_14617
n_14618
n_14619
n_14620
n_14621
n_14622
n_14623
n_14626
n_14627
n_14628
n_14629
n_1463
n_14631
n_14632
n_14633
n_14634
n_14636
n_14637
n_14638
n_14639
n_14640
n_14641
n_14643
n_14644
n_14646
n_14647
n_14648
n_14649
n_1465
n_14650
n_14651
n_14652
n_14653
n_14654
n_14655
n_14656
n_14657
n_14659
n_14660
n_14661
n_14663
n_14664
n_14665
n_14666
n_14667
n_14669
n_1467
n_14670
n_14671
n_14672
n_14673
n_14674
n_14675
n_14676
n_14678
n_14679
n_1468
n_14680
n_14681
n_14682
n_14683
n_14685
n_14686
n_14687
n_1469
n_14690
n_14693
n_14694
n_14695
n_14696
n_14697
n_14698
n_1470
n_14700
n_14701
n_14702
n_14703
n_14705
n_14706
n_14709
n_1471
n_14710
n_14711
n_14713
n_14715
n_14717
n_14719
n_1472
n_14721
n_14722
n_14723
n_14724
n_14725
n_14726
n_14727
n_14728
n_14731
n_14733
n_14734
n_14736
n_14738
n_1474
n_14740
n_14741
n_14743
n_14744
n_14746
n_14747
n_14748
n_14749
n_1475
n_14750
n_14751
n_14753
n_14754
n_14755
n_14756
n_14757
n_14759
n_1476
n_14760
n_14762
n_14763
n_14764
n_14766
n_14767
n_14768
n_14769
n_14772
n_14773
n_14775
n_14776
n_14777
n_14778
n_1478
n_14781
n_14783
n_14784
n_14786
n_14789
n_1479
n_14790
n_14791
n_14792
n_14793
n_14794
n_14796
n_14797
n_14798
n_14799
n_148
n_1480
n_14800
n_14802
n_14803
n_14804
n_14805
n_14806
n_14807
n_14808
n_1481
n_14810
n_14811
n_14812
n_14813
n_14814
n_14815
n_14816
n_14817
n_14818
n_14819
n_1482
n_14821
n_14822
n_14824
n_14825
n_14826
n_14828
n_14829
n_1483
n_14830
n_14832
n_14833
n_14834
n_14836
n_14837
n_14838
n_14839
n_1484
n_14840
n_14841
n_14842
n_14844
n_14845
n_14846
n_14847
n_14848
n_1485
n_14850
n_14851
n_14852
n_14853
n_14854
n_14855
n_14859
n_1486
n_14860
n_14861
n_14862
n_14864
n_14865
n_14866
n_14867
n_14869
n_14871
n_14873
n_14875
n_14877
n_14879
n_1488
n_14880
n_14881
n_14883
n_14884
n_14885
n_14887
n_14888
n_14889
n_14890
n_14891
n_14892
n_14894
n_14895
n_14896
n_14897
n_14898
n_14899
n_14900
n_14901
n_14902
n_14903
n_14904
n_14905
n_14906
n_14907
n_14908
n_14909
n_14910
n_14914
n_14916
n_14920
n_14921
n_14922
n_14923
n_14924
n_14930
n_14932
n_14933
n_1495
n_14956
n_14962
n_14963
n_14965
n_14967
n_1497
n_14971
n_14981
n_14987
n_1499
n_15
n_150
n_15001
n_1501
n_15014
n_1502
n_1503
n_15030
n_1504
n_15055
n_15065
n_1507
n_1508
n_1509
n_1510
n_15114
n_15115
n_15117
n_1512
n_15125
n_1513
n_15142
n_15188
n_1519
n_15190
n_15191
n_15204
n_15210
n_15217
n_1522
n_1523
n_15231
n_1524
n_15249
n_15260
n_15261
n_15275
n_15276
n_15291
n_15292
n_15295
n_15302
n_15313
n_1532
n_15324
n_15325
n_1533
n_15330
n_15331
n_15347
n_1535
n_15365
n_1537
n_15370
n_15371
n_15372
n_15373
n_15376
n_15377
n_15385
n_15388
n_15389
n_15390
n_15397
n_15403
n_15405
n_15407
n_1541
n_15438
n_15440
n_15441
n_15442
n_15444
n_15445
n_15446
n_1545
n_15453
n_15454
n_15456
n_15457
n_15458
n_1546
n_15467
n_15474
n_1548
n_1549
n_1551
n_15512
n_15513
n_15514
n_15515
n_15516
n_15517
n_15518
n_1552
n_15527
n_15528
n_15529
n_1553
n_15533
n_15534
n_15537
n_15538
n_15539
n_1554
n_15540
n_15549
n_1555
n_15551
n_15558
n_15565
n_15567
n_15568
n_1557
n_15576
n_1558
n_15587
n_1559
n_15592
n_15594
n_15596
n_15598
n_156
n_15601
n_15602
n_15604
n_15605
n_15607
n_1561
n_15611
n_15621
n_15625
n_15626
n_1563
n_15638
n_1564
n_15645
n_1565
n_1566
n_1567
n_15677
n_15680
n_15689
n_1569
n_15697
n_1570
n_1572
n_15726
n_15729
n_1573
n_15735
n_15736
n_15737
n_15738
n_15739
n_1574
n_15744
n_15746
n_15754
n_15755
n_15756
n_15757
n_15758
n_15759
n_15760
n_15761
n_15762
n_15763
n_15766
n_15768
n_15769
n_1577
n_15770
n_1578
n_15788
n_1579
n_15805
n_15808
n_1581
n_1582
n_15823
n_15824
n_15825
n_1583
n_1584
n_15841
n_15842
n_1585
n_15854
n_15856
n_15859
n_1586
n_1590
n_15908
n_15909
n_15910
n_15911
n_15914
n_15915
n_15916
n_15917
n_15918
n_15919
n_1592
n_15920
n_15921
n_15922
n_15923
n_15924
n_15927
n_15928
n_15929
n_1593
n_15931
n_15932
n_15935
n_15936
n_15937
n_15938
n_15939
n_1594
n_15940
n_15941
n_15942
n_1595
n_15958
n_15959
n_1596
n_15960
n_1597
n_15981
n_15988
n_1599
n_15994
n_15998
n_15999
n_160
n_1600
n_16000
n_16001
n_16002
n_16003
n_1601
n_16015
n_16016
n_16021
n_16027
n_1603
n_16030
n_16033
n_16034
n_16036
n_16046
n_16047
n_16048
n_16049
n_16052
n_1606
n_16066
n_1607
n_16070
n_16071
n_16075
n_16076
n_16089
n_1609
n_1610
n_16101
n_16102
n_16103
n_16105
n_1611
n_1612
n_1613
n_16131
n_1614
n_16150
n_16151
n_16152
n_16153
n_16154
n_16156
n_16158
n_16159
n_16160
n_16161
n_16162
n_16163
n_16164
n_16165
n_16166
n_16167
n_16168
n_16169
n_16170
n_16171
n_16172
n_16173
n_16175
n_16176
n_16181
n_16183
n_1619
n_16205
n_16206
n_16208
n_16209
n_1621
n_16210
n_16211
n_16212
n_16213
n_16224
n_1623
n_1624
n_16242
n_16243
n_16244
n_16247
n_16248
n_16249
n_1625
n_16250
n_16251
n_16252
n_16253
n_16254
n_1626
n_16262
n_16263
n_16264
n_16265
n_16268
n_16271
n_16273
n_16275
n_1628
n_16280
n_16284
n_16285
n_16286
n_16287
n_16288
n_16289
n_1629
n_16290
n_16291
n_16293
n_16297
n_16298
n_16299
n_1630
n_16300
n_16301
n_16303
n_16305
n_16306
n_16307
n_16310
n_16311
n_1632
n_16322
n_16325
n_16326
n_16327
n_1633
n_16331
n_16332
n_16338
n_1634
n_1635
n_16350
n_16351
n_16352
n_16354
n_16358
n_1636
n_16364
n_16368
n_16369
n_16370
n_16387
n_16388
n_16389
n_1639
n_16390
n_16391
n_16392
n_16393
n_16394
n_16395
n_16396
n_1640
n_16405
n_16408
n_16409
n_1641
n_16410
n_16411
n_16412
n_16413
n_1642
n_16424
n_16425
n_16427
n_16428
n_1643
n_16430
n_16431
n_16433
n_16434
n_16435
n_16436
n_16438
n_1644
n_16441
n_16442
n_16444
n_16451
n_16452
n_16456
n_1646
n_16460
n_16461
n_16462
n_1647
n_16474
n_16475
n_1648
n_16485
n_16486
n_16487
n_1649
n_16497
n_16499
n_1650
n_16500
n_16501
n_16503
n_16504
n_16506
n_16507
n_16508
n_16511
n_16512
n_16513
n_16516
n_16517
n_16518
n_16519
n_1652
n_16520
n_16521
n_16523
n_16524
n_1653
n_16533
n_16534
n_16535
n_16536
n_16538
n_1654
n_16541
n_16543
n_16544
n_16547
n_1655
n_16550
n_16553
n_16554
n_1656
n_16560
n_16564
n_16565
n_16566
n_1657
n_16572
n_16573
n_16574
n_16575
n_16576
n_16577
n_16578
n_16581
n_16582
n_16583
n_16584
n_16587
n_16591
n_16592
n_16594
n_16595
n_16598
n_16599
n_16601
n_16602
n_16603
n_16604
n_16605
n_16610
n_16612
n_16613
n_16614
n_16615
n_1662
n_16621
n_16622
n_16623
n_16626
n_16627
n_16628
n_16629
n_1663
n_16630
n_16631
n_16635
n_16637
n_1664
n_16657
n_1666
n_1667
n_1668
n_16685
n_1669
n_16690
n_16695
n_16696
n_16698
n_16720
n_1673
n_16735
n_16738
n_1674
n_16748
n_1675
n_16763
n_1677
n_16779
n_1678
n_1679
n_16791
n_16798
n_168
n_1680
n_1681
n_16810
n_16816
n_16818
n_1683
n_16834
n_16835
n_1684
n_16840
n_16841
n_16848
n_16849
n_16855
n_1686
n_16860
n_16864
n_16867
n_16871
n_16876
n_16888
n_1689
n_16891
n_169
n_1690
n_16904
n_16906
n_16914
n_16916
n_1692
n_1693
n_16934
n_16936
n_1694
n_16940
n_16942
n_16945
n_16949
n_1695
n_1696
n_16963
n_16964
n_16966
n_1697
n_16970
n_16974
n_16975
n_16976
n_16977
n_1698
n_16980
n_16981
n_16982
n_16984
n_16985
n_16986
n_16987
n_1699
n_16992
n_17
n_1700
n_1701
n_17013
n_17016
n_17017
n_17018
n_17019
n_17020
n_17021
n_17025
n_17027
n_17028
n_17029
n_17030
n_17034
n_17037
n_17038
n_17039
n_1704
n_17040
n_17041
n_17042
n_17043
n_17044
n_17045
n_17046
n_17047
n_17048
n_17049
n_17050
n_17051
n_1708
n_1709
n_1717
n_1719
n_1722
n_1724
n_1737
n_1739
n_1740
n_1742
n_1746
n_1748
n_1750
n_1752
n_1754
n_1755
n_1756
n_1758
n_1759
n_177
n_1774
n_1777
n_1779
n_1781
n_1782
n_1783
n_1784
n_1785
n_1786
n_1787
n_1788
n_1789
n_1790
n_1791
n_1793
n_1794
n_1795
n_1798
n_1799
n_18
n_1802
n_1803
n_1804
n_1805
n_1808
n_1809
n_1812
n_1813
n_1815
n_1816
n_1817
n_1819
n_1823
n_1824
n_1825
n_1826
n_1827
n_1828
n_1829
n_1830
n_1831
n_1832
n_1834
n_1835
n_1836
n_1837
n_1844
n_1845
n_1846
n_1847
n_1848
n_1851
n_1853
n_1854
n_1856
n_1857
n_1858
n_1859
n_1863
n_1864
n_1867
n_1868
n_1870
n_1871
n_1873
n_1874
n_1876
n_1877
n_1881
n_1882
n_1884
n_1885
n_1886
n_1887
n_1888
n_1889
n_1890
n_1891
n_1892
n_1894
n_1897
n_1899
n_1900
n_1902
n_1903
n_1904
n_1905
n_1907
n_1908
n_1909
n_191
n_1910
n_1911
n_1913
n_1914
n_1915
n_1916
n_1917
n_1918
n_1919
n_1920
n_1921
n_1922
n_1924
n_1926
n_1927
n_1928
n_1930
n_1931
n_1933
n_1934
n_1935
n_1937
n_1938
n_1939
n_1941
n_1942
n_1943
n_1944
n_1946
n_1948
n_1949
n_1950
n_1951
n_1952
n_1954
n_1956
n_1961
n_1963
n_1965
n_1966
n_1967
n_1968
n_1969
n_1970
n_1971
n_1972
n_1973
n_1976
n_1979
n_1981
n_1989
n_1990
n_1995
n_1996
n_1998
n_1999
n_2
n_200
n_2000
n_2001
n_2002
n_2004
n_2005
n_2006
n_2007
n_2008
n_2009
n_2010
n_2011
n_2012
n_2013
n_2015
n_2016
n_2017
n_2018
n_2019
n_202
n_2022
n_2023
n_2024
n_2027
n_2028
n_2031
n_2032
n_2033
n_2035
n_2036
n_2037
n_2038
n_204
n_2040
n_2041
n_2042
n_2044
n_2047
n_2048
n_2049
n_2051
n_2052
n_2053
n_2055
n_2057
n_2058
n_2059
n_2060
n_2065
n_2066
n_2067
n_2068
n_2069
n_207
n_2070
n_2071
n_2072
n_2075
n_2078
n_2079
n_2080
n_2084
n_2086
n_2087
n_2092
n_2093
n_2094
n_2100
n_2101
n_2102
n_2103
n_2104
n_2105
n_2106
n_2108
n_2110
n_2111
n_2113
n_2114
n_2115
n_2117
n_2119
n_2120
n_2121
n_2122
n_2125
n_2126
n_2127
n_2129
n_2131
n_2134
n_2135
n_2136
n_2137
n_2138
n_2146
n_2150
n_2151
n_2153
n_2154
n_2155
n_2156
n_2160
n_2161
n_2162
n_2163
n_2164
n_2165
n_2166
n_2168
n_2170
n_2171
n_2172
n_2173
n_2174
n_2175
n_2177
n_2178
n_2179
n_218
n_2180
n_2182
n_2183
n_2185
n_2186
n_2187
n_2188
n_2190
n_2191
n_2193
n_2194
n_2195
n_2196
n_2197
n_2198
n_2199
n_22
n_2201
n_2202
n_2204
n_2206
n_2207
n_2208
n_2209
n_221
n_2210
n_2211
n_2212
n_2213
n_2214
n_2215
n_2219
n_2223
n_2225
n_2226
n_2227
n_2228
n_2229
n_2230
n_2231
n_2232
n_2233
n_2235
n_2236
n_2237
n_2238
n_224
n_2241
n_2242
n_2243
n_2244
n_2245
n_2246
n_2247
n_2248
n_2250
n_2251
n_2253
n_2255
n_2256
n_2257
n_2258
n_2259
n_226
n_2260
n_2261
n_2263
n_2264
n_2266
n_2267
n_2269
n_2271
n_2272
n_2273
n_2274
n_2275
n_2276
n_228
n_2280
n_2281
n_2284
n_2285
n_2289
n_229
n_2291
n_2292
n_2293
n_2295
n_2297
n_2298
n_2299
n_23
n_230
n_2300
n_2301
n_2302
n_2304
n_2305
n_2306
n_2308
n_2311
n_2313
n_2314
n_2315
n_2316
n_2319
n_232
n_2326
n_2327
n_2329
n_233
n_2331
n_2337
n_2339
n_234
n_2341
n_2343
n_2344
n_2345
n_2347
n_2349
n_235
n_2350
n_2352
n_2353
n_2356
n_2358
n_2359
n_236
n_2361
n_2362
n_2363
n_2364
n_2366
n_2367
n_2369
n_2371
n_2373
n_2375
n_2376
n_2377
n_2380
n_2381
n_2387
n_2388
n_2389
n_239
n_2390
n_2392
n_2395
n_2396
n_2397
n_2398
n_2399
n_2400
n_2401
n_2403
n_2404
n_2405
n_2406
n_2407
n_2409
n_2410
n_2411
n_2412
n_2414
n_2415
n_2416
n_2418
n_2419
n_2420
n_2421
n_2423
n_2424
n_2426
n_2427
n_2428
n_2429
n_243
n_2430
n_2431
n_2432
n_2433
n_2434
n_2435
n_2436
n_2437
n_2438
n_2439
n_2440
n_2441
n_2442
n_2445
n_2446
n_2447
n_2449
n_2451
n_2453
n_2456
n_2457
n_2458
n_2459
n_2460
n_2461
n_2462
n_2463
n_2464
n_2468
n_2469
n_2473
n_2475
n_2476
n_2477
n_2478
n_2479
n_2482
n_2483
n_2485
n_2486
n_2487
n_2488
n_249
n_2491
n_2492
n_2493
n_2494
n_2496
n_2497
n_2498
n_2499
n_2500
n_2501
n_2502
n_2503
n_2504
n_2505
n_2508
n_2509
n_251
n_2510
n_2512
n_2513
n_2514
n_2515
n_2516
n_2517
n_2518
n_2519
n_2520
n_2521
n_2522
n_2524
n_2526
n_2527
n_2528
n_2530
n_2531
n_2533
n_2536
n_2537
n_2539
n_2540
n_2541
n_2542
n_2543
n_2544
n_2545
n_2547
n_255
n_2552
n_2553
n_2555
n_2556
n_2558
n_2560
n_2562
n_2564
n_2566
n_2567
n_2568
n_2569
n_257
n_2570
n_2571
n_2572
n_2573
n_2574
n_2575
n_2577
n_2579
n_2580
n_2581
n_2582
n_2584
n_2585
n_2587
n_2588
n_2590
n_2592
n_2594
n_2595
n_2596
n_2597
n_2598
n_2599
n_26
n_2601
n_2602
n_2603
n_2604
n_2605
n_2606
n_2608
n_2609
n_261
n_2610
n_2612
n_2613
n_2615
n_2616
n_2619
n_262
n_2620
n_2622
n_2623
n_2624
n_2625
n_2627
n_2629
n_263
n_2630
n_2631
n_2632
n_2633
n_2634
n_2635
n_2636
n_2637
n_2638
n_2639
n_264
n_2640
n_2641
n_2643
n_2645
n_2646
n_2648
n_2649
n_265
n_2651
n_2652
n_2654
n_2655
n_2657
n_2659
n_2661
n_2663
n_2664
n_2665
n_2666
n_2670
n_2671
n_2673
n_2674
n_2675
n_2676
n_2677
n_2678
n_2679
n_268
n_2680
n_2681
n_2682
n_2684
n_2685
n_2687
n_2691
n_2692
n_2693
n_2694
n_2695
n_2696
n_2697
n_2698
n_2699
n_2700
n_2701
n_2702
n_2704
n_2705
n_2706
n_2707
n_2708
n_2709
n_271
n_2710
n_2711
n_2712
n_2713
n_2714
n_2715
n_2716
n_2717
n_2719
n_272
n_2720
n_2721
n_2722
n_2723
n_2725
n_2727
n_2728
n_2729
n_2730
n_2732
n_2734
n_2735
n_2738
n_2739
n_2740
n_2742
n_2744
n_2745
n_2748
n_2750
n_2751
n_2752
n_2753
n_2754
n_2755
n_2756
n_2757
n_276
n_2761
n_2762
n_2763
n_2764
n_2767
n_2768
n_2769
n_277
n_2770
n_2774
n_2776
n_2777
n_2778
n_2779
n_278
n_2780
n_2781
n_2782
n_2783
n_2784
n_2785
n_2786
n_2787
n_2788
n_2789
n_279
n_2790
n_2792
n_2793
n_2795
n_2799
n_2804
n_2806
n_2807
n_2809
n_2812
n_2813
n_2814
n_2815
n_282
n_2820
n_2822
n_2825
n_2828
n_2829
n_2831
n_2835
n_2838
n_2841
n_2842
n_2844
n_285
n_2850
n_2851
n_2852
n_2854
n_2855
n_2858
n_2860
n_2864
n_2866
n_2867
n_2868
n_2869
n_287
n_2870
n_2871
n_2872
n_2873
n_2874
n_2876
n_2877
n_2878
n_288
n_2888
n_2897
n_2902
n_2904
n_2907
n_2909
n_2910
n_2911
n_2914
n_2915
n_2916
n_2917
n_2918
n_2919
n_292
n_2920
n_2921
n_2922
n_2924
n_2925
n_2929
n_2931
n_2932
n_2933
n_2934
n_2935
n_2937
n_2938
n_2939
n_2940
n_2941
n_2942
n_2943
n_2947
n_2948
n_2949
n_295
n_2950
n_2952
n_2953
n_2954
n_2955
n_2956
n_2957
n_2958
n_2959
n_2960
n_2961
n_2962
n_2964
n_2966
n_2967
n_2968
n_297
n_2970
n_2971
n_2972
n_2979
n_298
n_2980
n_2981
n_2982
n_2983
n_2986
n_2987
n_2988
n_2989
n_2990
n_2991
n_2992
n_2993
n_2995
n_2997
n_2998
n_2999
n_300
n_3000
n_3001
n_3004
n_3005
n_3006
n_3007
n_3008
n_3013
n_3014
n_3015
n_3016
n_3017
n_3018
n_3019
n_3020
n_3021
n_3022
n_3024
n_3025
n_3026
n_3027
n_3028
n_303
n_3030
n_3031
n_3032
n_3033
n_3034
n_3036
n_304
n_3044
n_3046
n_3048
n_3049
n_305
n_3050
n_3052
n_3054
n_3055
n_3057
n_3058
n_306
n_3061
n_3064
n_3066
n_3068
n_3071
n_3072
n_3076
n_3077
n_3080
n_3083
n_3084
n_3087
n_3089
n_3090
n_3107
n_3108
n_3110
n_3111
n_3112
n_3113
n_3114
n_3115
n_3116
n_3118
n_3119
n_3120
n_3123
n_3125
n_313
n_3130
n_3131
n_3132
n_3133
n_3134
n_3135
n_3136
n_3137
n_3138
n_3139
n_3140
n_3141
n_3142
n_3147
n_3148
n_3151
n_3152
n_3153
n_3154
n_3156
n_3157
n_3158
n_3159
n_3160
n_3162
n_3164
n_3166
n_3167
n_3168
n_3169
n_317
n_3170
n_3171
n_3172
n_3173
n_3174
n_3175
n_3178
n_3179
n_3185
n_3189
n_319
n_3190
n_3191
n_3192
n_3193
n_3194
n_3195
n_3196
n_3197
n_3198
n_3199
n_320
n_3200
n_3201
n_3202
n_3203
n_3204
n_3205
n_3206
n_3207
n_321
n_3210
n_3211
n_3212
n_3213
n_3214
n_3215
n_3216
n_3217
n_3219
n_3220
n_3221
n_3222
n_3223
n_3224
n_3226
n_3228
n_3229
n_323
n_3231
n_3233
n_3237
n_3238
n_324
n_3241
n_3246
n_3248
n_325
n_3250
n_3251
n_3252
n_3253
n_3254
n_3255
n_3256
n_3257
n_3258
n_3259
n_3261
n_3262
n_3265
n_3266
n_3267
n_3268
n_3269
n_3271
n_3273
n_3274
n_3275
n_3276
n_3277
n_3278
n_3279
n_3280
n_3281
n_3282
n_3283
n_3284
n_3285
n_3286
n_3289
n_329
n_3290
n_3293
n_3294
n_3295
n_3296
n_3297
n_3298
n_3301
n_3302
n_3304
n_3305
n_3306
n_331
n_3310
n_3313
n_3314
n_3315
n_3316
n_3317
n_3318
n_3319
n_3320
n_3321
n_3323
n_3324
n_3325
n_3326
n_3327
n_333
n_3330
n_3331
n_3332
n_3333
n_3334
n_3335
n_3337
n_3338
n_3339
n_3340
n_3341
n_3342
n_3344
n_3345
n_3346
n_3347
n_3348
n_3349
n_335
n_3350
n_3351
n_3352
n_3353
n_3354
n_3355
n_3356
n_3357
n_3358
n_3359
n_3360
n_3361
n_3363
n_3364
n_3365
n_3366
n_3367
n_3368
n_3370
n_3371
n_3372
n_3373
n_3374
n_3375
n_3376
n_3377
n_3381
n_3384
n_3385
n_3386
n_3387
n_3388
n_3389
n_3390
n_3391
n_3392
n_3393
n_3395
n_3399
n_34
n_340
n_3402
n_3407
n_3409
n_341
n_3410
n_3413
n_3414
n_3415
n_3416
n_3417
n_3419
n_342
n_3420
n_3421
n_3422
n_3423
n_3425
n_3426
n_3427
n_3428
n_343
n_3432
n_3436
n_3438
n_3440
n_3445
n_3448
n_3449
n_345
n_3452
n_3453
n_3454
n_3456
n_3457
n_3458
n_3459
n_3460
n_3461
n_3463
n_3464
n_3465
n_3466
n_3467
n_3468
n_3469
n_3470
n_3471
n_3472
n_3474
n_3475
n_3476
n_3477
n_3478
n_3479
n_3480
n_3481
n_3482
n_3483
n_3484
n_3485
n_3486
n_3487
n_3488
n_3489
n_349
n_3490
n_3491
n_3492
n_3493
n_3494
n_3496
n_3497
n_3498
n_3499
n_350
n_3501
n_3502
n_3503
n_3504
n_3506
n_3507
n_3508
n_3509
n_351
n_3510
n_3511
n_3515
n_3517
n_3519
n_3523
n_3524
n_3527
n_3528
n_3530
n_3531
n_3533
n_3537
n_3538
n_3539
n_3542
n_3543
n_3544
n_3546
n_3547
n_3549
n_355
n_3550
n_3552
n_3553
n_3555
n_3556
n_3557
n_3558
n_3560
n_3563
n_3564
n_3565
n_3570
n_3572
n_3573
n_3574
n_3577
n_3579
n_358
n_3580
n_3582
n_3583
n_3584
n_3586
n_3588
n_3589
n_3590
n_3591
n_3592
n_3593
n_3596
n_3597
n_3598
n_3599
n_36
n_360
n_3600
n_3601
n_3602
n_3607
n_3608
n_3609
n_3610
n_3613
n_3615
n_3616
n_3617
n_3618
n_362
n_3621
n_3622
n_3623
n_3624
n_3625
n_3626
n_3627
n_3628
n_3629
n_3630
n_3634
n_3638
n_364
n_3641
n_3642
n_3643
n_3644
n_3645
n_3647
n_3649
n_3651
n_3652
n_3654
n_3655
n_3659
n_366
n_3660
n_3661
n_3662
n_3664
n_3665
n_3666
n_3667
n_3670
n_3671
n_3674
n_3676
n_3677
n_3678
n_3680
n_3681
n_3683
n_3684
n_3694
n_3695
n_3696
n_3697
n_3699
n_370
n_3700
n_3701
n_3702
n_3703
n_3704
n_3705
n_3706
n_3707
n_3710
n_3711
n_3713
n_3714
n_3715
n_3717
n_3719
n_372
n_3720
n_3721
n_3722
n_3724
n_3725
n_3727
n_3729
n_373
n_3730
n_3731
n_3732
n_3737
n_3739
n_374
n_3741
n_3744
n_3745
n_3746
n_3747
n_3749
n_375
n_3750
n_3751
n_3752
n_3755
n_3757
n_376
n_3761
n_3762
n_3763
n_3764
n_3765
n_3769
n_377
n_3770
n_3771
n_3772
n_3773
n_3774
n_3776
n_3777
n_3778
n_3779
n_3780
n_3781
n_3783
n_3784
n_3785
n_3786
n_3788
n_3789
n_3791
n_3792
n_3793
n_3794
n_3795
n_3796
n_3797
n_3798
n_38
n_3805
n_3806
n_3807
n_3808
n_3809
n_3810
n_3811
n_3813
n_3816
n_3817
n_3819
n_382
n_3820
n_3822
n_3823
n_3824
n_3825
n_3827
n_3829
n_3831
n_3832
n_3833
n_3834
n_3835
n_3839
n_384
n_3844
n_3845
n_3847
n_3849
n_385
n_3851
n_3852
n_3853
n_3854
n_3856
n_386
n_3860
n_3862
n_3863
n_3864
n_3865
n_3866
n_3868
n_3870
n_3872
n_3874
n_3875
n_3876
n_3877
n_3879
n_3880
n_3882
n_3883
n_3884
n_3885
n_3887
n_3889
n_389
n_3891
n_3893
n_3895
n_3897
n_390
n_3900
n_3901
n_3904
n_3905
n_3906
n_3909
n_391
n_3914
n_3917
n_3918
n_392
n_3921
n_3922
n_3923
n_3926
n_3927
n_3928
n_3929
n_3933
n_3935
n_3937
n_3938
n_3940
n_3941
n_3944
n_3945
n_3947
n_3950
n_3953
n_3954
n_3955
n_3956
n_3958
n_3959
n_396
n_3960
n_3961
n_3965
n_3967
n_3968
n_3969
n_397
n_3973
n_3976
n_3977
n_3978
n_3979
n_3980
n_3981
n_3982
n_3983
n_3984
n_3987
n_3988
n_3989
n_3990
n_3991
n_3993
n_3994
n_3995
n_3996
n_3997
n_40
n_4000
n_4002
n_4003
n_4007
n_4008
n_4009
n_401
n_4010
n_4012
n_4013
n_4016
n_4017
n_4019
n_4021
n_4022
n_4023
n_4024
n_4029
n_403
n_4030
n_4031
n_4032
n_4035
n_4036
n_4037
n_4038
n_4039
n_404
n_4041
n_4043
n_4045
n_4047
n_4048
n_4049
n_405
n_4050
n_4051
n_4053
n_4054
n_4056
n_4058
n_4060
n_4061
n_4065
n_407
n_4071
n_4073
n_4074
n_4076
n_4077
n_4078
n_408
n_4080
n_4084
n_4085
n_4086
n_409
n_4090
n_4092
n_4093
n_4095
n_4098
n_4100
n_4105
n_4106
n_4107
n_4108
n_4109
n_411
n_4111
n_4112
n_4113
n_4114
n_4115
n_4119
n_412
n_4123
n_413
n_4130
n_4131
n_4132
n_4134
n_4135
n_4136
n_4137
n_4138
n_4140
n_4142
n_4143
n_4149
n_415
n_4151
n_4152
n_4153
n_4154
n_4157
n_4158
n_4159
n_4160
n_4161
n_4162
n_4163
n_4165
n_4168
n_4169
n_4170
n_4171
n_4172
n_4177
n_4178
n_418
n_4188
n_419
n_4190
n_4191
n_4192
n_4193
n_4195
n_4196
n_4197
n_4198
n_4199
n_42
n_420
n_4200
n_4201
n_4203
n_4204
n_4205
n_4206
n_4207
n_4208
n_4209
n_4210
n_4211
n_4212
n_4213
n_4214
n_4216
n_4217
n_4218
n_4219
n_4223
n_4228
n_4229
n_4231
n_4233
n_4234
n_4235
n_4238
n_424
n_4241
n_4242
n_4243
n_4244
n_4248
n_425
n_4250
n_4254
n_4255
n_4258
n_4260
n_4262
n_4263
n_4265
n_4271
n_4273
n_4274
n_4276
n_4277
n_4278
n_4279
n_4282
n_4284
n_4285
n_4286
n_4287
n_4290
n_4292
n_4293
n_4295
n_4296
n_4297
n_4298
n_430
n_4303
n_4304
n_4305
n_4308
n_4314
n_4318
n_432
n_4320
n_4327
n_4328
n_4329
n_433
n_4330
n_4331
n_4334
n_4336
n_4339
n_434
n_4340
n_4341
n_4345
n_4346
n_4347
n_4348
n_435
n_4350
n_4351
n_4352
n_4353
n_4354
n_4357
n_4361
n_4365
n_4366
n_4369
n_4372
n_4373
n_4374
n_4376
n_4378
n_4379
n_438
n_4380
n_4381
n_4382
n_4383
n_4385
n_4386
n_4388
n_4389
n_4390
n_440
n_4401
n_4402
n_4406
n_4407
n_4413
n_4414
n_4415
n_4417
n_4419
n_4420
n_4421
n_4427
n_4431
n_4433
n_4434
n_4437
n_4438
n_4439
n_4442
n_4444
n_4445
n_4446
n_4447
n_4450
n_4452
n_4454
n_4457
n_4458
n_4459
n_4460
n_4465
n_4467
n_4468
n_4470
n_4471
n_4473
n_4474
n_4475
n_4476
n_4478
n_4479
n_4480
n_4482
n_4484
n_4485
n_4487
n_4488
n_4489
n_4493
n_4494
n_4496
n_4498
n_4501
n_4504
n_4506
n_4507
n_4509
n_4512
n_4513
n_4514
n_4515
n_4516
n_4517
n_4518
n_4520
n_4521
n_4522
n_4523
n_4524
n_4525
n_4527
n_4528
n_4532
n_4533
n_4534
n_4535
n_4536
n_4537
n_4592
n_4593
n_4594
n_4595
n_46
n_4601
n_4603
n_4605
n_4607
n_4610
n_4612
n_4614
n_4616
n_4619
n_4621
n_4623
n_4625
n_4627
n_4628
n_4629
n_4630
n_4631
n_4632
n_4633
n_4634
n_4635
n_4636
n_4637
n_4638
n_4639
n_4642
n_4644
n_4645
n_4647
n_4649
n_4658
n_4662
n_4666
n_4667
n_4668
n_4669
n_4671
n_4672
n_4674
n_4675
n_4676
n_4677
n_4678
n_4680
n_4681
n_4686
n_4687
n_4688
n_4690
n_4692
n_4693
n_4694
n_4696
n_4697
n_4698
n_4700
n_4701
n_4702
n_4704
n_4705
n_4706
n_4707
n_4708
n_471
n_4710
n_4711
n_4712
n_4713
n_4714
n_4715
n_4716
n_4717
n_4718
n_4720
n_4721
n_4722
n_4723
n_4724
n_4725
n_4726
n_4727
n_4728
n_4729
n_4730
n_4732
n_4733
n_4734
n_4736
n_4737
n_4739
n_4740
n_4741
n_4743
n_4744
n_4746
n_4747
n_4748
n_4749
n_4750
n_4751
n_4752
n_4753
n_4754
n_4755
n_4756
n_4757
n_4758
n_4759
n_4760
n_4761
n_4762
n_4763
n_4764
n_4765
n_4766
n_4767
n_4768
n_4769
n_4770
n_4771
n_4772
n_4773
n_4774
n_4775
n_4776
n_4777
n_4778
n_4779
n_4781
n_4782
n_4783
n_4784
n_4785
n_4786
n_4787
n_4795
n_4796
n_4797
n_4798
n_4799
n_4802
n_4803
n_4806
n_4812
n_4814
n_4815
n_4816
n_4818
n_4819
n_4820
n_4822
n_4823
n_4828
n_4830
n_4831
n_4832
n_4833
n_4834
n_4835
n_4836
n_4837
n_4838
n_4840
n_4841
n_4842
n_4843
n_4844
n_4845
n_4846
n_4847
n_4848
n_4853
n_4854
n_4856
n_4862
n_4863
n_4864
n_4866
n_4867
n_4868
n_4869
n_4871
n_4872
n_4873
n_4874
n_4875
n_4877
n_4878
n_4879
n_4880
n_4881
n_4882
n_4884
n_4885
n_4886
n_4887
n_4888
n_4889
n_4890
n_4891
n_4893
n_4894
n_4895
n_4896
n_4897
n_4900
n_4901
n_4902
n_4903
n_4904
n_4906
n_4909
n_4911
n_4912
n_4913
n_4914
n_4917
n_4918
n_4920
n_4922
n_4924
n_4926
n_4928
n_4930
n_4932
n_4934
n_4936
n_4939
n_4943
n_4945
n_4949
n_4951
n_4955
n_4963
n_497
n_4973
n_4975
n_4980
n_4982
n_4984
n_4986
n_4991
n_4996
n_4999
n_5003
n_5009
n_5012
n_5018
n_5021
n_5023
n_5025
n_5027
n_5029
n_5036
n_5038
n_504
n_5042
n_5044
n_5048
n_5052
n_5054
n_5058
n_5060
n_5066
n_5071
n_5074
n_5078
n_5082
n_5088
n_5092
n_5094
n_5096
n_5100
n_5102
n_5104
n_5112
n_5116
n_5118
n_512
n_5122
n_5124
n_513
n_5130
n_5136
n_5138
n_5140
n_5143
n_5149
n_5151
n_5163
n_5168
n_5170
n_5176
n_5179
n_518
n_5185
n_5188
n_519
n_5192
n_5198
n_520
n_5207
n_521
n_5210
n_5212
n_5216
n_5218
n_522
n_5223
n_5225
n_5227
n_523
n_5230
n_5237
n_524
n_5244
n_5246
n_525
n_5251
n_5253
n_5255
n_5260
n_527
n_5272
n_5277
n_5279
n_528
n_529
n_5293
n_5296
n_530
n_5300
n_5303
n_5305
n_531
n_5313
n_5315
n_5318
n_5323
n_5325
n_5327
n_533
n_5335
n_534
n_5342
n_5349
n_5351
n_5361
n_5368
n_5371
n_5373
n_5376
n_5378
n_5383
n_5386
n_5388
n_539
n_5391
n_5393
n_5399
n_540
n_5402
n_5406
n_541
n_5412
n_5414
n_5416
n_5418
n_5421
n_5424
n_5427
n_5435
n_5438
n_5441
n_5444
n_5446
n_5450
n_5452
n_5454
n_5456
n_5458
n_546
n_5461
n_5465
n_547
n_5474
n_5478
n_5481
n_5483
n_5486
n_5489
n_549
n_5491
n_5493
n_550
n_5501
n_5503
n_5505
n_5507
n_5509
n_551
n_5513
n_5515
n_5517
n_5521
n_5526
n_5528
n_5534
n_5537
n_554
n_5541
n_5545
n_5546
n_5547
n_5548
n_5549
n_5553
n_5556
n_5557
n_5558
n_5559
n_5561
n_5563
n_5565
n_5567
n_5568
n_5569
n_5571
n_5573
n_5574
n_5575
n_5577
n_5578
n_558
n_5580
n_5582
n_5583
n_5587
n_5588
n_5589
n_559
n_5592
n_5594
n_5595
n_5597
n_5600
n_5603
n_5614
n_5616
n_5618
n_5619
n_5620
n_5622
n_5623
n_5625
n_5626
n_5627
n_5628
n_5632
n_5633
n_5639
n_564
n_5640
n_5641
n_5644
n_5645
n_5648
n_5649
n_565
n_5651
n_5652
n_5655
n_5657
n_5658
n_566
n_5660
n_5663
n_5666
n_5668
n_567
n_5670
n_5672
n_5673
n_5675
n_5676
n_5678
n_5679
n_568
n_5681
n_5682
n_5684
n_5686
n_5688
n_5689
n_5691
n_5694
n_5696
n_5699
n_57
n_5702
n_5703
n_5705
n_5708
n_5709
n_5710
n_5712
n_5717
n_5722
n_5723
n_5725
n_5729
n_573
n_5731
n_5732
n_5733
n_5736
n_574
n_5740
n_5742
n_5743
n_5744
n_5745
n_5747
n_5749
n_5750
n_5751
n_5752
n_5753
n_5754
n_5755
n_5757
n_5763
n_5766
n_5768
n_5769
n_5770
n_5774
n_5776
n_5778
n_5780
n_5784
n_5788
n_5790
n_5798
n_580
n_5802
n_5806
n_581
n_5810
n_582
n_5822
n_583
n_5838
n_584
n_5840
n_5842
n_5844
n_5848
n_585
n_5850
n_5854
n_5858
n_586
n_5860
n_5862
n_5866
n_587
n_5876
n_588
n_5880
n_5882
n_589
n_5896
n_5898
n_5904
n_5906
n_5920
n_5922
n_593
n_5930
n_5934
n_5936
n_594
n_5940
n_5944
n_595
n_5954
n_5958
n_596
n_5960
n_5962
n_5964
n_5967
n_597
n_5971
n_5975
n_5979
n_598
n_5981
n_5983
n_5989
n_599
n_5999
n_6
n_600
n_6001
n_6005
n_6007
n_601
n_6011
n_6013
n_6015
n_6019
n_602
n_6023
n_6027
n_6029
n_6033
n_604
n_6040
n_6041
n_6043
n_6045
n_6049
n_6051
n_6054
n_606
n_6060
n_6063
n_6067
n_6069
n_607
n_6071
n_6073
n_6077
n_6079
n_609
n_6091
n_6095
n_6099
n_61
n_610
n_6101
n_6103
n_6105
n_6107
n_6109
n_611
n_6111
n_6115
n_612
n_6125
n_6132
n_6135
n_6136
n_6138
n_614
n_6142
n_6146
n_615
n_6152
n_6158
n_616
n_6162
n_6168
n_617
n_6173
n_6177
n_6181
n_6186
n_6189
n_6191
n_6193
n_6195
n_6199
n_620
n_6200
n_6201
n_6206
n_6211
n_622
n_6221
n_6223
n_6226
n_6228
n_6230
n_6231
n_6232
n_6240
n_6246
n_6249
n_625
n_6254
n_6257
n_6259
n_626
n_6261
n_6266
n_6268
n_627
n_6271
n_6273
n_6276
n_6278
n_6281
n_6284
n_6286
n_6287
n_629
n_6292
n_6295
n_6297
n_6298
n_6303
n_6313
n_6319
n_6325
n_6327
n_6329
n_6337
n_6340
n_6342
n_6344
n_6347
n_6348
n_6350
n_6361
n_6364
n_6366
n_6369
n_6371
n_6376
n_6382
n_6386
n_6388
n_639
n_6390
n_6391
n_640
n_6400
n_6402
n_6405
n_641
n_6410
n_6413
n_6415
n_642
n_6420
n_6423
n_6425
n_6427
n_643
n_6431
n_6435
n_6436
n_6443
n_6446
n_6448
n_645
n_6453
n_6456
n_646
n_6461
n_6465
n_6468
n_6475
n_6477
n_648
n_6483
n_6488
n_649
n_6495
n_6498
n_65
n_650
n_6504
n_6509
n_6512
n_6516
n_6518
n_652
n_6521
n_653
n_6530
n_6534
n_6538
n_654
n_6543
n_655
n_6550
n_6553
n_6554
n_6556
n_656
n_6561
n_6567
n_657
n_6572
n_6575
n_6578
n_6582
n_6587
n_659
n_6594
n_6596
n_6603
n_6605
n_6613
n_6615
n_662
n_6620
n_6621
n_6623
n_6626
n_6629
n_663
n_6634
n_6639
n_664
n_6644
n_6645
n_6651
n_6654
n_6659
n_666
n_6662
n_6665
n_6674
n_668
n_6682
n_6684
n_669
n_6693
n_6697
n_67
n_670
n_6703
n_6707
n_6709
n_6716
n_6718
n_6726
n_6729
n_6735
n_6738
n_674
n_6745
n_6749
n_675
n_6752
n_6757
n_6768
n_677
n_6772
n_6776
n_678
n_6783
n_6785
n_6788
n_6791
n_6793
n_6799
n_6801
n_6804
n_6809
n_681
n_6812
n_6816
n_6819
n_6824
n_6826
n_6828
n_6830
n_6835
n_6840
n_6842
n_6849
n_6853
n_6855
n_6861
n_6867
n_6868
n_6869
n_6871
n_6872
n_6885
n_6886
n_6887
n_689
n_6892
n_6895
n_6897
n_6898
n_6902
n_6903
n_691
n_6917
n_692
n_6920
n_6926
n_6932
n_6934
n_6935
n_6937
n_6941
n_6943
n_6944
n_6946
n_695
n_6951
n_6953
n_6956
n_696
n_6971
n_6980
n_6983
n_6986
n_6988
n_6989
n_6991
n_6996
n_700
n_7003
n_7004
n_7005
n_7006
n_7007
n_7010
n_7012
n_7013
n_7015
n_7016
n_7018
n_7019
n_7027
n_7029
n_7030
n_7032
n_7033
n_7034
n_7038
n_7039
n_7040
n_7043
n_7044
n_7045
n_7046
n_7047
n_7048
n_705
n_7050
n_7051
n_7052
n_7053
n_7054
n_7056
n_7057
n_706
n_7060
n_7061
n_7062
n_7063
n_7065
n_7067
n_7070
n_7071
n_7072
n_7073
n_7074
n_7075
n_7078
n_708
n_7080
n_7081
n_7082
n_7083
n_7084
n_7085
n_7086
n_7087
n_7088
n_7089
n_709
n_7091
n_7092
n_7095
n_7096
n_7108
n_711
n_7110
n_7112
n_7114
n_7115
n_7117
n_7119
n_7121
n_7122
n_7123
n_7125
n_7126
n_7128
n_713
n_7130
n_7132
n_7134
n_7135
n_7136
n_7137
n_7139
n_7141
n_7143
n_7145
n_7147
n_7149
n_7151
n_7153
n_7155
n_7157
n_7159
n_7161
n_7163
n_7165
n_7168
n_7171
n_7174
n_7177
n_7180
n_7182
n_7185
n_7187
n_7189
n_7191
n_7193
n_7195
n_7197
n_7200
n_7203
n_7205
n_7207
n_7209
n_721
n_7211
n_7213
n_7214
n_7215
n_7216
n_7217
n_7218
n_7219
n_7223
n_7224
n_7225
n_7226
n_7227
n_7231
n_7233
n_7234
n_7235
n_7239
n_7240
n_7241
n_7242
n_7244
n_7249
n_7252
n_7253
n_7256
n_7257
n_7259
n_7260
n_7262
n_7264
n_7265
n_7266
n_7267
n_7268
n_7269
n_727
n_7270
n_7272
n_7273
n_7274
n_7275
n_7276
n_7277
n_7278
n_7279
n_7281
n_7282
n_7283
n_7287
n_7288
n_7289
n_729
n_7291
n_7293
n_7294
n_7295
n_7296
n_7297
n_7298
n_730
n_7308
n_7309
n_731
n_7310
n_7311
n_7312
n_7313
n_7316
n_7317
n_7320
n_7321
n_7322
n_7324
n_7325
n_7326
n_7327
n_7329
n_733
n_7330
n_7334
n_7335
n_7337
n_7338
n_7339
n_734
n_7341
n_7344
n_7350
n_736
n_7362
n_7368
n_7369
n_737
n_7371
n_7373
n_7375
n_7377
n_7379
n_738
n_7383
n_7385
n_7386
n_7387
n_7388
n_739
n_7390
n_7396
n_7397
n_7399
n_74
n_740
n_7401
n_7405
n_7406
n_7408
n_741
n_7410
n_7411
n_7412
n_7415
n_7417
n_7418
n_742
n_7420
n_7421
n_7422
n_7423
n_7424
n_7425
n_7426
n_7427
n_7428
n_743
n_7430
n_7431
n_7432
n_7433
n_7437
n_7438
n_744
n_7440
n_7442
n_7443
n_7444
n_7445
n_7446
n_7447
n_7448
n_7449
n_745
n_7450
n_7451
n_7454
n_746
n_7464
n_7466
n_747
n_7470
n_7476
n_7478
n_7479
n_748
n_7480
n_7481
n_7482
n_7485
n_7487
n_7488
n_7489
n_7490
n_7492
n_7493
n_7495
n_7497
n_7498
n_7499
n_7500
n_7504
n_7505
n_7507
n_7508
n_7509
n_7510
n_7511
n_7512
n_7513
n_7514
n_7516
n_7517
n_7518
n_7519
n_7521
n_7522
n_7523
n_7524
n_7525
n_7527
n_7529
n_7530
n_7531
n_7532
n_7534
n_7535
n_7538
n_7540
n_7541
n_7547
n_7551
n_7552
n_7557
n_7558
n_7559
n_7560
n_7561
n_7562
n_7564
n_7565
n_7567
n_7569
n_7574
n_7575
n_7577
n_7578
n_7580
n_7582
n_7583
n_7586
n_7587
n_7588
n_7589
n_7591
n_7592
n_7593
n_7594
n_7596
n_7597
n_7598
n_76
n_7603
n_7608
n_7609
n_7614
n_7615
n_7616
n_7617
n_7618
n_7619
n_7620
n_7622
n_7624
n_7626
n_7627
n_7629
n_763
n_7631
n_7633
n_7635
n_7638
n_7639
n_7640
n_7642
n_7645
n_7647
n_7648
n_7649
n_7650
n_7651
n_7652
n_7653
n_7656
n_7657
n_7664
n_7665
n_7666
n_7667
n_7669
n_7671
n_7672
n_7673
n_7677
n_7679
n_7681
n_7683
n_7684
n_7685
n_7687
n_7689
n_7692
n_7694
n_7695
n_7697
n_7698
n_7699
n_7701
n_7702
n_7703
n_7704
n_7705
n_7706
n_7707
n_7708
n_7709
n_7710
n_7711
n_7712
n_7715
n_7716
n_7717
n_7720
n_7721
n_7722
n_7724
n_7725
n_7726
n_7729
n_7730
n_7731
n_7733
n_7734
n_7735
n_7737
n_7738
n_7739
n_7740
n_7744
n_7746
n_7747
n_7749
n_7750
n_7751
n_7752
n_7753
n_7754
n_7755
n_7756
n_7757
n_7759
n_7760
n_7761
n_7762
n_7766
n_7767
n_7768
n_7769
n_7771
n_7773
n_7774
n_7776
n_7777
n_7779
n_7780
n_7781
n_7782
n_7783
n_7785
n_7786
n_7787
n_7788
n_7789
n_779
n_7790
n_7791
n_7792
n_7795
n_7796
n_7797
n_7798
n_7799
n_7800
n_7801
n_7802
n_7803
n_7804
n_7805
n_7806
n_7807
n_7808
n_7809
n_7810
n_7811
n_7812
n_7813
n_7814
n_7815
n_7818
n_7821
n_7822
n_7823
n_7824
n_7826
n_7828
n_7830
n_7833
n_7835
n_7836
n_7838
n_7840
n_7842
n_7844
n_7845
n_7849
n_7851
n_7853
n_7859
n_7861
n_7863
n_7865
n_7867
n_7869
n_7873
n_7879
n_7881
n_7883
n_7889
n_7891
n_7893
n_7895
n_7897
n_7899
n_790
n_7901
n_7903
n_7905
n_7907
n_7909
n_7911
n_7915
n_7917
n_7919
n_7923
n_7925
n_7927
n_7931
n_7935
n_7937
n_7939
n_7945
n_7947
n_7949
n_7953
n_7955
n_7957
n_7959
n_7961
n_7963
n_7965
n_7967
n_7969
n_7971
n_7973
n_7975
n_7977
n_798
n_7981
n_7985
n_7989
n_7991
n_7993
n_7995
n_7997
n_8001
n_8005
n_8012
n_8014
n_8017
n_802
n_8021
n_8024
n_8027
n_8030
n_8032
n_8034
n_8036
n_8039
n_8041
n_8044
n_8047
n_8049
n_8052
n_8056
n_8059
n_8060
n_8068
n_8069
n_8071
n_8073
n_8076
n_8079
n_808
n_8082
n_8084
n_8087
n_8094
n_8097
n_8100
n_8107
n_8109
n_8111
n_8114
n_8116
n_8118
n_8119
n_812
n_8121
n_8123
n_8128
n_813
n_8132
n_8135
n_8137
n_8139
n_8140
n_8142
n_815
n_8150
n_8159
n_816
n_8161
n_8163
n_8168
n_817
n_8171
n_8173
n_8175
n_8176
n_8178
n_8180
n_8182
n_8184
n_8186
n_8189
n_819
n_8191
n_8193
n_8196
n_8200
n_8203
n_8205
n_8210
n_8213
n_8215
n_8220
n_8229
n_8232
n_8239
n_824
n_8241
n_8244
n_8248
n_8251
n_8253
n_8255
n_8258
n_826
n_8260
n_8262
n_8264
n_8267
n_8269
n_8271
n_8272
n_8274
n_8277
n_8281
n_8283
n_8285
n_829
n_8291
n_8293
n_8295
n_8299
n_83
n_8304
n_8307
n_8309
n_8316
n_8319
n_8321
n_8323
n_8325
n_8327
n_8329
n_8331
n_8333
n_8335
n_8337
n_8339
n_834
n_8341
n_8344
n_8346
n_8349
n_835
n_8351
n_8353
n_8355
n_8358
n_836
n_8360
n_8364
n_8366
n_8368
n_837
n_8371
n_8373
n_838
n_8382
n_8384
n_839
n_8391
n_8393
n_8395
n_8397
n_84
n_840
n_8400
n_8402
n_8404
n_8406
n_8407
n_8409
n_841
n_8411
n_8413
n_8415
n_8417
n_8419
n_842
n_8421
n_8423
n_8426
n_843
n_8430
n_8431
n_8433
n_8434
n_8436
n_8437
n_8438
n_8439
n_844
n_8440
n_8441
n_8442
n_8444
n_8446
n_8447
n_8448
n_8449
n_845
n_8450
n_8451
n_8452
n_8455
n_8456
n_8457
n_8458
n_8459
n_846
n_8460
n_8461
n_8462
n_8463
n_8464
n_8465
n_8466
n_8467
n_8468
n_8469
n_847
n_8470
n_8472
n_8476
n_8478
n_848
n_8480
n_8481
n_8483
n_8486
n_8487
n_8488
n_8489
n_849
n_8492
n_8493
n_8494
n_8495
n_8496
n_8498
n_850
n_8500
n_8501
n_8502
n_8503
n_8504
n_8505
n_8506
n_8509
n_851
n_8511
n_8512
n_8513
n_8514
n_8515
n_8516
n_8517
n_8518
n_8519
n_852
n_8520
n_8521
n_8522
n_8523
n_8524
n_8526
n_8527
n_853
n_8535
n_8538
n_8540
n_8541
n_8542
n_8547
n_8548
n_855
n_8551
n_8558
n_856
n_8561
n_8564
n_8565
n_8566
n_8567
n_8568
n_8569
n_857
n_8570
n_8571
n_8572
n_8573
n_8576
n_8579
n_858
n_8580
n_8582
n_8585
n_8588
n_8589
n_859
n_8590
n_8591
n_8595
n_860
n_8601
n_8602
n_8603
n_8604
n_8605
n_8606
n_8607
n_861
n_8616
n_8617
n_8618
n_8619
n_862
n_8620
n_8621
n_8622
n_8623
n_8624
n_8625
n_8626
n_8627
n_8628
n_8629
n_863
n_8630
n_8631
n_8632
n_8633
n_8634
n_8635
n_8636
n_8637
n_8638
n_864
n_8640
n_8641
n_8642
n_8643
n_8644
n_8645
n_8646
n_8647
n_865
n_8652
n_8653
n_8657
n_8658
n_8659
n_866
n_8660
n_8664
n_8668
n_8669
n_867
n_8672
n_8674
n_8678
n_868
n_8682
n_8688
n_869
n_8692
n_8693
n_8694
n_8695
n_8697
n_8699
n_870
n_8701
n_8703
n_8705
n_8707
n_8708
n_8709
n_871
n_8711
n_8713
n_8714
n_8716
n_8717
n_872
n_8721
n_8724
n_8725
n_8726
n_8727
n_8728
n_873
n_8730
n_8731
n_8732
n_8733
n_8734
n_8736
n_8738
n_874
n_8740
n_8741
n_8742
n_8743
n_8744
n_8745
n_8746
n_8747
n_8748
n_875
n_8751
n_8756
n_8757
n_8759
n_876
n_8765
n_877
n_878
n_8784
n_879
n_8790
n_8794
n_8795
n_880
n_8800
n_8801
n_881
n_8818
n_8819
n_882
n_8820
n_883
n_8831
n_8832
n_8833
n_8834
n_8835
n_8837
n_8838
n_884
n_8840
n_8841
n_8842
n_8843
n_8846
n_8847
n_8848
n_8849
n_885
n_8850
n_8851
n_8852
n_8853
n_8854
n_8855
n_8856
n_8857
n_8859
n_886
n_8860
n_8863
n_8864
n_8866
n_8867
n_887
n_8871
n_8872
n_8874
n_8875
n_8876
n_8877
n_8879
n_888
n_8884
n_889
n_8892
n_8896
n_8897
n_8898
n_8899
n_890
n_8908
n_891
n_8910
n_8917
n_8919
n_892
n_8920
n_8921
n_8924
n_8926
n_8927
n_8928
n_893
n_8932
n_8934
n_8939
n_894
n_8940
n_8941
n_8944
n_8946
n_8949
n_895
n_8950
n_8951
n_8953
n_8954
n_8955
n_8960
n_8962
n_8963
n_8964
n_8970
n_8971
n_8973
n_8977
n_8979
n_898
n_8981
n_8983
n_8986
n_899
n_8992
n_8993
n_8994
n_8996
n_900
n_9001
n_9002
n_9003
n_9004
n_9007
n_9008
n_9009
n_901
n_9010
n_9011
n_9012
n_9013
n_9014
n_9015
n_9016
n_9017
n_9018
n_9019
n_902
n_9020
n_9022
n_9023
n_9025
n_9026
n_9027
n_9028
n_903
n_9032
n_9033
n_9034
n_9035
n_904
n_9041
n_9044
n_9045
n_9046
n_9047
n_9048
n_9049
n_905
n_9051
n_9054
n_9056
n_9057
n_9058
n_9059
n_906
n_9060
n_9061
n_9062
n_9063
n_9064
n_9066
n_9067
n_9068
n_9069
n_907
n_9070
n_9071
n_9072
n_9074
n_9075
n_9076
n_9077
n_9078
n_908
n_9080
n_9081
n_9086
n_9088
n_909
n_9090
n_9093
n_9094
n_9096
n_9097
n_9098
n_9099
n_910
n_9100
n_9102
n_9103
n_9104
n_9105
n_9106
n_9107
n_9108
n_911
n_9110
n_9111
n_9112
n_9113
n_9115
n_9116
n_9117
n_9118
n_9119
n_912
n_9120
n_9121
n_9122
n_9123
n_9124
n_9125
n_9126
n_9127
n_9129
n_913
n_9131
n_9133
n_9134
n_9137
n_914
n_9141
n_9142
n_9143
n_9144
n_9145
n_9146
n_915
n_9152
n_9153
n_9154
n_9155
n_9157
n_916
n_9160
n_9163
n_9168
n_917
n_9170
n_9171
n_9172
n_9173
n_9174
n_9175
n_9176
n_9177
n_9178
n_9179
n_918
n_9180
n_9181
n_9182
n_9183
n_9184
n_9185
n_9187
n_9188
n_9189
n_919
n_9192
n_9197
n_9198
n_920
n_9200
n_9202
n_9203
n_9204
n_9206
n_9209
n_921
n_9215
n_9216
n_9218
n_9219
n_922
n_9220
n_9221
n_9222
n_9223
n_9224
n_9226
n_9228
n_9229
n_923
n_9232
n_9233
n_9234
n_9235
n_9236
n_9237
n_9238
n_9239
n_924
n_9241
n_9256
n_926
n_9260
n_9265
n_9269
n_927
n_9271
n_9272
n_9274
n_9276
n_9277
n_928
n_9284
n_9285
n_9286
n_9287
n_929
n_9290
n_9293
n_9294
n_9295
n_9296
n_9297
n_9298
n_9299
n_930
n_9301
n_9307
n_9309
n_931
n_9311
n_9312
n_9315
n_9319
n_9320
n_9321
n_9322
n_9329
n_9330
n_9331
n_9332
n_9334
n_9335
n_9340
n_9341
n_9342
n_9343
n_9345
n_9346
n_9348
n_9350
n_9353
n_9355
n_9358
n_9361
n_9363
n_9366
n_9368
n_937
n_9371
n_9372
n_9374
n_9377
n_9379
n_938
n_9381
n_9383
n_9385
n_9387
n_9389
n_939
n_9391
n_9393
n_9396
n_9398
n_940
n_9400
n_9402
n_9404
n_9406
n_9407
n_9408
n_941
n_9410
n_9411
n_9412
n_9414
n_9416
n_9418
n_9419
n_9420
n_9421
n_9423
n_9426
n_9427
n_9428
n_943
n_9430
n_9431
n_9435
n_9436
n_9437
n_9438
n_9439
n_944
n_9440
n_9442
n_9443
n_9444
n_9445
n_9446
n_9447
n_9448
n_9449
n_945
n_9450
n_9451
n_9453
n_9454
n_9455
n_9456
n_9457
n_9459
n_946
n_9460
n_9461
n_9463
n_9464
n_9465
n_9467
n_9468
n_9469
n_947
n_9470
n_9471
n_9472
n_9473
n_9474
n_9475
n_9476
n_9477
n_9478
n_948
n_9481
n_9485
n_9486
n_9487
n_9488
n_9489
n_949
n_9490
n_9492
n_9493
n_9494
n_9495
n_9496
n_9497
n_9498
n_9499
n_95
n_950
n_9500
n_9502
n_9504
n_9505
n_9506
n_9507
n_9508
n_951
n_9510
n_9512
n_9513
n_9514
n_9515
n_9516
n_9517
n_9518
n_9519
n_952
n_9520
n_9521
n_9522
n_9523
n_9524
n_9525
n_9526
n_9527
n_9528
n_9529
n_9531
n_9532
n_9534
n_9537
n_9538
n_9539
n_9540
n_9541
n_9542
n_9543
n_9544
n_9545
n_9546
n_9547
n_9548
n_955
n_9550
n_9551
n_9552
n_9553
n_9554
n_9555
n_9557
n_9558
n_9559
n_956
n_9560
n_9561
n_9565
n_9568
n_9569
n_957
n_9570
n_9571
n_9572
n_9573
n_9575
n_9576
n_9578
n_9579
n_958
n_9583
n_9584
n_9586
n_9588
n_959
n_9590
n_9591
n_9592
n_9593
n_9594
n_9596
n_9598
n_960
n_9600
n_9602
n_9604
n_9605
n_9607
n_961
n_9610
n_9613
n_9615
n_9617
n_9619
n_9621
n_9624
n_9625
n_9626
n_963
n_9631
n_9633
n_9635
n_9637
n_9639
n_964
n_9640
n_9642
n_9645
n_9648
n_9649
n_965
n_9651
n_9653
n_9657
n_9659
n_9660
n_9663
n_9665
n_9666
n_9667
n_9668
n_9669
n_9671
n_9673
n_9674
n_9676
n_9677
n_9682
n_9683
n_9684
n_9686
n_9687
n_9689
n_969
n_9690
n_9691
n_9692
n_9693
n_9694
n_9696
n_9697
n_9700
n_9701
n_9703
n_9705
n_9706
n_9707
n_9708
n_9709
n_971
n_9710
n_9711
n_9712
n_9713
n_9714
n_9715
n_9717
n_9718
n_9719
n_9721
n_9722
n_9723
n_9724
n_9725
n_9726
n_9728
n_973
n_9731
n_9732
n_9733
n_9734
n_9735
n_9737
n_9738
n_974
n_9740
n_9741
n_9744
n_9747
n_9752
n_9753
n_9754
n_9756
n_9757
n_9759
n_976
n_9761
n_9765
n_9776
n_9779
n_978
n_9781
n_9785
n_9789
n_9790
n_9791
n_9793
n_9794
n_9796
n_9798
n_980
n_9800
n_9802
n_9804
n_9807
n_9811
n_9814
n_9816
n_9818
n_982
n_9822
n_9823
n_9825
n_9826
n_9827
n_9828
n_983
n_9830
n_9831
n_9832
n_9833
n_9834
n_9835
n_9836
n_9837
n_9838
n_9839
n_9840
n_9841
n_9842
n_9843
n_9844
n_9845
n_9846
n_9847
n_9849
n_9850
n_9851
n_9852
n_9853
n_9854
n_9855
n_9856
n_9857
n_9858
n_9859
n_9860
n_9861
n_9862
n_9863
n_9864
n_9865
n_9868
n_987
n_9872
n_9874
n_9875
n_9876
n_9877
n_9878
n_9879
n_988
n_9880
n_9881
n_9882
n_9883
n_9884
n_9885
n_9886
n_9888
n_9889
n_9890
n_9891
n_9892
n_9894
n_9895
n_9896
n_9897
n_9898
n_9899
n_990
n_9901
n_9902
n_9903
n_9904
n_9906
n_9908
n_9912
n_9914
n_9916
n_992
n_9926
n_9928
n_993
n_9931
n_9932
n_994
n_9941
n_9942
n_9947
n_9950
n_9953
n_996
n_9968
n_9971
n_9976
n_9979
n_998
n_9988
n_999
n_9992
n_9997
output_backup_devsel_out_reg_Q
output_backup_par_en_out_reg_Q
output_backup_par_out_reg_Q
output_backup_serr_en_out_reg_Q
output_backup_stop_out_reg_Q
output_backup_tar_ad_en_out_reg_Q
output_backup_trdy_out_reg_Q
parchk_pci_ad_out_in
parchk_pci_ad_out_in_1168
parchk_pci_ad_out_in_1169
parchk_pci_ad_out_in_1170
parchk_pci_ad_out_in_1171
parchk_pci_ad_out_in_1172
parchk_pci_ad_out_in_1173
parchk_pci_ad_out_in_1174
parchk_pci_ad_out_in_1175
parchk_pci_ad_out_in_1177
parchk_pci_ad_out_in_1178
parchk_pci_ad_out_in_1179
parchk_pci_ad_out_in_1180
parchk_pci_ad_out_in_1181
parchk_pci_ad_out_in_1182
parchk_pci_ad_out_in_1183
parchk_pci_ad_out_in_1184
parchk_pci_ad_out_in_1185
parchk_pci_ad_out_in_1186
parchk_pci_ad_out_in_1187
parchk_pci_ad_out_in_1188
parchk_pci_ad_out_in_1191
parchk_pci_ad_out_in_1192
parchk_pci_ad_out_in_1193
parchk_pci_ad_out_in_1194
parchk_pci_ad_out_in_1197
parchk_pci_ad_reg_in
parchk_pci_ad_reg_in_1205
parchk_pci_ad_reg_in_1206
parchk_pci_ad_reg_in_1207
parchk_pci_ad_reg_in_1208
parchk_pci_ad_reg_in_1209
parchk_pci_ad_reg_in_1210
parchk_pci_ad_reg_in_1211
parchk_pci_ad_reg_in_1212
parchk_pci_ad_reg_in_1213
parchk_pci_ad_reg_in_1214
parchk_pci_ad_reg_in_1215
parchk_pci_ad_reg_in_1216
parchk_pci_ad_reg_in_1217
parchk_pci_ad_reg_in_1218
parchk_pci_ad_reg_in_1219
parchk_pci_ad_reg_in_1220
parchk_pci_ad_reg_in_1221
parchk_pci_ad_reg_in_1222
parchk_pci_ad_reg_in_1223
parchk_pci_ad_reg_in_1224
parchk_pci_ad_reg_in_1225
parchk_pci_ad_reg_in_1226
parchk_pci_ad_reg_in_1227
parchk_pci_ad_reg_in_1228
parchk_pci_ad_reg_in_1229
parchk_pci_ad_reg_in_1230
parchk_pci_ad_reg_in_1231
parchk_pci_ad_reg_in_1232
parchk_pci_ad_reg_in_1233
parchk_pci_ad_reg_in_1235
parchk_pci_cbe_en_in
parchk_pci_cbe_out_in
parchk_pci_cbe_out_in_1202
parchk_pci_cbe_out_in_1203
parchk_pci_cbe_out_in_1204
parchk_pci_cbe_reg_in
parchk_pci_cbe_reg_in_1236
parchk_pci_cbe_reg_in_1237
parchk_pci_cbe_reg_in_1238
parchk_pci_frame_reg_in
parchk_pci_par_en_in
parchk_pci_serr_en_in
parchk_pci_serr_out_in
parchk_pci_trdy_en_in
parity_checker_check_for_serr_on_second
parity_checker_check_for_serr_on_second_reg_Q
parity_checker_frame_and_irdy_en_prev
parity_checker_frame_and_irdy_en_prev_prev
parity_checker_frame_dec2
parity_checker_master_perr_report
parity_checker_master_perr_report_reg_Q
pci_inti_conf_int_in
pci_target_unit_del_sync_addr_in
pci_target_unit_del_sync_addr_in_205
pci_target_unit_del_sync_addr_in_206
pci_target_unit_del_sync_addr_in_207
pci_target_unit_del_sync_addr_in_208
pci_target_unit_del_sync_addr_in_209
pci_target_unit_del_sync_addr_in_210
pci_target_unit_del_sync_addr_in_212
pci_target_unit_del_sync_addr_in_213
pci_target_unit_del_sync_addr_in_214
pci_target_unit_del_sync_addr_in_217
pci_target_unit_del_sync_addr_in_218
pci_target_unit_del_sync_addr_in_219
pci_target_unit_del_sync_addr_in_220
pci_target_unit_del_sync_addr_in_221
pci_target_unit_del_sync_addr_in_222
pci_target_unit_del_sync_addr_in_223
pci_target_unit_del_sync_addr_in_224
pci_target_unit_del_sync_addr_in_225
pci_target_unit_del_sync_addr_in_226
pci_target_unit_del_sync_addr_in_227
pci_target_unit_del_sync_addr_in_228
pci_target_unit_del_sync_addr_in_230
pci_target_unit_del_sync_addr_in_231
pci_target_unit_del_sync_addr_in_232
pci_target_unit_del_sync_addr_in_233
pci_target_unit_del_sync_addr_in_234
pci_target_unit_del_sync_bc_in
pci_target_unit_del_sync_bc_in_201
pci_target_unit_del_sync_bc_in_202
pci_target_unit_del_sync_bc_in_203
pci_target_unit_del_sync_be_out_reg_0__Q
pci_target_unit_del_sync_be_out_reg_1__Q
pci_target_unit_del_sync_be_out_reg_2__Q
pci_target_unit_del_sync_be_out_reg_3__Q
pci_target_unit_del_sync_comp_cycle_count_0_
pci_target_unit_del_sync_comp_cycle_count_10_
pci_target_unit_del_sync_comp_cycle_count_11_
pci_target_unit_del_sync_comp_cycle_count_12_
pci_target_unit_del_sync_comp_cycle_count_13_
pci_target_unit_del_sync_comp_cycle_count_14_
pci_target_unit_del_sync_comp_cycle_count_15_
pci_target_unit_del_sync_comp_cycle_count_1_
pci_target_unit_del_sync_comp_cycle_count_2_
pci_target_unit_del_sync_comp_cycle_count_3_
pci_target_unit_del_sync_comp_cycle_count_4_
pci_target_unit_del_sync_comp_cycle_count_5_
pci_target_unit_del_sync_comp_cycle_count_6_
pci_target_unit_del_sync_comp_cycle_count_7_
pci_target_unit_del_sync_comp_cycle_count_8_
pci_target_unit_del_sync_comp_cycle_count_9_
pci_target_unit_del_sync_comp_cycle_count_reg_16__Q
pci_target_unit_del_sync_comp_done_reg_clr
pci_target_unit_del_sync_comp_done_reg_clr_reg_Q
pci_target_unit_del_sync_comp_done_reg_main
pci_target_unit_del_sync_comp_done_reg_main_reg_Q
pci_target_unit_del_sync_comp_in
pci_target_unit_del_sync_comp_rty_exp_clr
pci_target_unit_del_sync_comp_rty_exp_clr_reg_Q
pci_target_unit_del_sync_comp_rty_exp_reg
pci_target_unit_del_sync_req_comp_pending
pci_target_unit_del_sync_req_comp_pending_sample
pci_target_unit_del_sync_req_comp_pending_sample_reg_Q
pci_target_unit_del_sync_req_done_reg
pci_target_unit_del_sync_req_rty_exp_clr
pci_target_unit_del_sync_req_rty_exp_clr_reg_Q
pci_target_unit_del_sync_req_rty_exp_reg
pci_target_unit_del_sync_req_sync_sync_data_out_reg_0__Q
pci_target_unit_del_sync_sync_comp_done
pci_target_unit_del_sync_sync_comp_req_pending
pci_target_unit_del_sync_sync_comp_rty_exp_clr
pci_target_unit_del_sync_sync_req_comp_pending
pci_target_unit_del_sync_sync_req_rty_exp
pci_target_unit_fifos_inGreyCount_0_
pci_target_unit_fifos_inGreyCount_reg_0__Q
pci_target_unit_fifos_inGreyCount_reg_1__Q
pci_target_unit_fifos_outGreyCount_0_
pci_target_unit_fifos_outGreyCount_reg_0__Q
pci_target_unit_fifos_outGreyCount_reg_1__Q
pci_target_unit_fifos_pcir_control_in_192
pci_target_unit_fifos_pcir_data_in
pci_target_unit_fifos_pcir_data_in_158
pci_target_unit_fifos_pcir_data_in_159
pci_target_unit_fifos_pcir_data_in_160
pci_target_unit_fifos_pcir_data_in_161
pci_target_unit_fifos_pcir_data_in_162
pci_target_unit_fifos_pcir_data_in_163
pci_target_unit_fifos_pcir_data_in_164
pci_target_unit_fifos_pcir_data_in_165
pci_target_unit_fifos_pcir_data_in_166
pci_target_unit_fifos_pcir_data_in_167
pci_target_unit_fifos_pcir_data_in_168
pci_target_unit_fifos_pcir_data_in_169
pci_target_unit_fifos_pcir_data_in_170
pci_target_unit_fifos_pcir_data_in_171
pci_target_unit_fifos_pcir_data_in_172
pci_target_unit_fifos_pcir_data_in_173
pci_target_unit_fifos_pcir_data_in_174
pci_target_unit_fifos_pcir_data_in_175
pci_target_unit_fifos_pcir_data_in_176
pci_target_unit_fifos_pcir_data_in_177
pci_target_unit_fifos_pcir_data_in_178
pci_target_unit_fifos_pcir_data_in_179
pci_target_unit_fifos_pcir_data_in_180
pci_target_unit_fifos_pcir_data_in_181
pci_target_unit_fifos_pcir_data_in_182
pci_target_unit_fifos_pcir_data_in_183
pci_target_unit_fifos_pcir_data_in_184
pci_target_unit_fifos_pcir_data_in_185
pci_target_unit_fifos_pcir_data_in_186
pci_target_unit_fifos_pcir_data_in_187
pci_target_unit_fifos_pcir_data_in_188
pci_target_unit_fifos_pcir_fifo_ctrl_raddr_1_
pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_1_
pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_2_
pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg_0__Q
pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg_2__Q
pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg_0__Q
pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg_1__Q
pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg_2__Q
pci_target_unit_fifos_pcir_fifo_ctrl_rclk_sync_wgrey_addr
pci_target_unit_fifos_pcir_fifo_ctrl_rclk_sync_wgrey_addr_39
pci_target_unit_fifos_pcir_fifo_ctrl_rclk_sync_wgrey_addr_40
pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_0_
pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_1_
pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_2_
pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg_0__Q
pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg_1__Q
pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg_2__Q
pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_0_
pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_1_
pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_2_
pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg_0__Q
pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg_1__Q
pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg_2__Q
pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_0_
pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_1_
pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_2_
pci_target_unit_fifos_pcir_fifo_ctrl_wclk_sync_rgrey_addr
pci_target_unit_fifos_pcir_fifo_ctrl_wclk_sync_rgrey_addr_100
pci_target_unit_fifos_pcir_fifo_ctrl_wclk_sync_rgrey_addr_101
pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg_0__Q
pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg_1__Q
pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg_2__Q
pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_0_
pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_1_
pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_2_
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__0__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__11__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__12__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__13__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__14__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__15__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__16__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__17__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__18__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__19__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__1__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__20__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__21__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__24__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__25__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__26__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__29__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__2__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__30__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__31__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__37__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__3__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__4__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__5__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__6__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__8__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__9__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__0__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__11__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__12__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__13__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__14__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__15__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__16__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__17__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__18__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__19__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__1__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__20__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__21__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__22__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__24__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__25__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__26__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__29__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__2__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__30__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__31__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__37__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__3__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__4__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__5__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__9__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__0__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__11__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__12__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__13__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__14__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__15__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__16__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__17__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__18__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__19__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__1__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__20__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__21__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__22__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__24__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__25__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__26__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__29__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__2__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__30__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__37__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__3__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__4__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__5__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__6__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__8__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__0__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__11__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__12__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__13__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__14__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__15__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__16__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__17__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__18__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__19__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__1__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__20__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__21__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__22__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__24__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__25__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__26__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__29__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__2__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__30__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__31__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__37__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__4__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__5__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__6__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__8__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__9__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__0__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__11__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__12__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__13__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__14__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__15__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__16__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__17__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__18__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__19__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__1__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__20__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__21__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__22__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__23__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__24__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__25__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__26__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__29__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__2__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__37__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__3__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__4__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__5__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__6__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__8__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__9__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__0__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__10__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__11__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__12__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__13__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__14__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__15__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__16__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__17__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__18__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__19__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__1__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__20__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__21__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__22__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__23__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__24__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__25__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__26__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__29__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__2__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__30__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__37__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__3__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__4__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__5__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__6__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__8__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__9__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__0__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__11__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__12__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__13__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__14__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__15__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__16__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__17__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__18__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__19__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__1__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__20__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__21__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__22__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__24__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__25__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__26__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__2__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__37__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__3__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__4__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__5__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__6__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__8__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__9__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__0__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__11__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__12__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__13__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__14__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__15__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__16__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__17__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__18__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__19__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__1__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__20__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__21__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__22__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__24__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__25__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__26__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__2__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__37__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__3__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__4__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__5__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__6__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__8__Q
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__9__Q
pci_target_unit_fifos_pcir_flush_in
pci_target_unit_fifos_pcir_wenable_in
pci_target_unit_fifos_pcir_whole_waddr
pci_target_unit_fifos_pcir_whole_waddr_94
pci_target_unit_fifos_pciw_addr_data_in
pci_target_unit_fifos_pciw_addr_data_in_121
pci_target_unit_fifos_pciw_addr_data_in_122
pci_target_unit_fifos_pciw_addr_data_in_123
pci_target_unit_fifos_pciw_addr_data_in_125
pci_target_unit_fifos_pciw_addr_data_in_126
pci_target_unit_fifos_pciw_addr_data_in_127
pci_target_unit_fifos_pciw_addr_data_in_128
pci_target_unit_fifos_pciw_addr_data_in_130
pci_target_unit_fifos_pciw_addr_data_in_131
pci_target_unit_fifos_pciw_addr_data_in_132
pci_target_unit_fifos_pciw_addr_data_in_133
pci_target_unit_fifos_pciw_addr_data_in_134
pci_target_unit_fifos_pciw_addr_data_in_135
pci_target_unit_fifos_pciw_addr_data_in_136
pci_target_unit_fifos_pciw_addr_data_in_137
pci_target_unit_fifos_pciw_addr_data_in_138
pci_target_unit_fifos_pciw_addr_data_in_139
pci_target_unit_fifos_pciw_addr_data_in_140
pci_target_unit_fifos_pciw_addr_data_in_141
pci_target_unit_fifos_pciw_addr_data_in_142
pci_target_unit_fifos_pciw_addr_data_in_143
pci_target_unit_fifos_pciw_addr_data_in_145
pci_target_unit_fifos_pciw_addr_data_in_146
pci_target_unit_fifos_pciw_addr_data_in_147
pci_target_unit_fifos_pciw_addr_data_in_148
pci_target_unit_fifos_pciw_addr_data_in_149
pci_target_unit_fifos_pciw_addr_data_in_150
pci_target_unit_fifos_pciw_addr_data_in_151
pci_target_unit_fifos_pciw_cbe_in
pci_target_unit_fifos_pciw_cbe_in_152
pci_target_unit_fifos_pciw_cbe_in_153
pci_target_unit_fifos_pciw_cbe_in_154
pci_target_unit_fifos_pciw_control_in
pci_target_unit_fifos_pciw_control_in_155
pci_target_unit_fifos_pciw_control_in_156
pci_target_unit_fifos_pciw_control_in_157
pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg_0__Q
pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg_1__Q
pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg_2__Q
pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg_0__Q
pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg_1__Q
pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg_2__Q
pci_target_unit_fifos_pciw_fifo_ctrl_rclk_sync_wgrey_addr
pci_target_unit_fifos_pciw_fifo_ctrl_rclk_sync_wgrey_addr_74
pci_target_unit_fifos_pciw_fifo_ctrl_rclk_sync_wgrey_addr_75
pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_0_
pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_1_
pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_2_
pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_0_
pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_1_
pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_2_
pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus1_reg_0__Q
pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus1_reg_1__Q
pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus1_reg_2__Q
pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus2_reg_0__Q
pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus2_reg_1__Q
pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus2_reg_2__Q
pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg_0__Q
pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg_1__Q
pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg_2__Q
pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_0_
pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_1_
pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_2_
pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_0_
pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_1_
pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_2_
pci_target_unit_fifos_pciw_fifo_ctrl_wclk_sync_rgrey_minus2
pci_target_unit_fifos_pciw_fifo_ctrl_wclk_sync_rgrey_minus_94
pci_target_unit_fifos_pciw_fifo_ctrl_wclk_sync_rgrey_minus_95
pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_0_
pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_1_
pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_2_
pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_0_
pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_1_
pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_2_
pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_0_
pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_1_
pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_2_
pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_0_
pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_1_
pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_2_
pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_37__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_0__153
pci_target_unit_fifos_pciw_fifo_storage_mem_1__192
pci_target_unit_fifos_pciw_fifo_storage_mem_2__231
pci_target_unit_fifos_pciw_fifo_storage_mem_3__270
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__10__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__11__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__13__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__14__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__16__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__17__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__20__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__22__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__23__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__25__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__26__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__28__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__29__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__2__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__30__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__32__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__33__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__34__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__36__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__37__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__38__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__39__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__3__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__8__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__0__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__10__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__11__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__13__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__17__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__1__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__20__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__22__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__23__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__25__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__26__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__28__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__29__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__2__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__30__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__32__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__33__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__34__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__35__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__36__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__37__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__38__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__39__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__3__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__6__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__8__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__0__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__10__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__11__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__14__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__15__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__17__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__18__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__20__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__22__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__23__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__25__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__26__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__29__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__2__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__30__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__31__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__32__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__33__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__34__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__35__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__36__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__37__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__38__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__39__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__3__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__6__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__8__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__0__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__10__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__11__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__14__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__15__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__17__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__18__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__20__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__22__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__23__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__25__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__26__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__27__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__29__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__2__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__30__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__31__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__32__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__33__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__34__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__36__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__37__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__38__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__39__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__3__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__5__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__8__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__10__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__12__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__15__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__17__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__18__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__21__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__22__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__23__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__25__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__26__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__28__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__29__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__2__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__30__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__32__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__33__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__34__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__35__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__36__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__37__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__38__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__39__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__3__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__5__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__6__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__8__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__0__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__10__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__12__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__14__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__17__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__18__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__20__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__21__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__22__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__23__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__25__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__28__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__29__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__2__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__30__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__32__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__33__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__34__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__35__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__36__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__37__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__38__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__39__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__3__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__5__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__6__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__8__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__0__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__10__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__13__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__15__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__17__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__18__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__21__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__22__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__23__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__25__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__26__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__29__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__2__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__30__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__31__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__32__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__33__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__34__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__35__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__36__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__37__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__38__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__39__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__3__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__5__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__6__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__8__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__10__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__12__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__13__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__15__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__17__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__18__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__20__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__21__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__23__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__25__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__26__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__27__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__29__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__2__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__30__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__31__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__32__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__33__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__34__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__35__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__36__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__37__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__38__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__39__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__3__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__6__Q
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__8__Q
pci_target_unit_fifos_pciw_inTransactionCount_0_
pci_target_unit_fifos_pciw_inTransactionCount_1_
pci_target_unit_fifos_pciw_inTransactionCount_reg_1__Q
pci_target_unit_fifos_pciw_outTransactionCount_1_
pci_target_unit_fifos_pciw_outTransactionCount_reg_0__Q
pci_target_unit_fifos_pciw_outTransactionCount_reg_1__Q
pci_target_unit_fifos_pciw_wenable_in
pci_target_unit_fifos_pciw_whole_waddr
pci_target_unit_fifos_pciw_whole_waddr_47
pci_target_unit_fifos_wb_clk_inGreyCount_0_
pci_target_unit_fifos_wb_clk_inGreyCount_1_
pci_target_unit_fifos_wb_clk_sync_inGreyCount
pci_target_unit_fifos_wb_clk_sync_inGreyCount_36
pci_target_unit_pci_target_if_async_reset_as_pcir_flush_async_reset_data_out_reg_Q
pci_target_unit_pci_target_if_keep_desconnect_wo_data_set
pci_target_unit_pci_target_if_norm_address_reg_0__Q
pci_target_unit_pci_target_if_norm_address_reg_2__Q
pci_target_unit_pci_target_if_norm_address_reg_3__Q
pci_target_unit_pci_target_if_norm_address_reg_4__Q
pci_target_unit_pci_target_if_norm_address_reg_5__Q
pci_target_unit_pci_target_if_norm_address_reg_6__Q
pci_target_unit_pci_target_if_norm_address_reg_7__Q
pci_target_unit_pci_target_if_norm_address_reg_9__Q
pci_target_unit_pci_target_if_norm_prf_en
pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_0__Q
pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_10__Q
pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_11__Q
pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_12__Q
pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_13__Q
pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_14__Q
pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_15__Q
pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_16__Q
pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_17__Q
pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_18__Q
pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_19__Q
pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_1__Q
pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_20__Q
pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_21__Q
pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_22__Q
pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_23__Q
pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_24__Q
pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_25__Q
pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_26__Q
pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_27__Q
pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_28__Q
pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_29__Q
pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_2__Q
pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_30__Q
pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_31__Q
pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_3__Q
pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_4__Q
pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_5__Q
pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_6__Q
pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_7__Q
pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_8__Q
pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_9__Q
pci_target_unit_pci_target_if_pciw_fifo_control_out_reg_0__Q
pci_target_unit_pci_target_if_same_read_reg
pci_target_unit_pci_target_sm_cnf_progress
pci_target_unit_pci_target_sm_n_2
pci_target_unit_pci_target_sm_n_3
pci_target_unit_pci_target_sm_rd_progress
pci_target_unit_pci_target_sm_read_completed_reg
pci_target_unit_pci_target_sm_read_completed_reg_reg_Q
pci_target_unit_pci_target_sm_same_read_reg
pci_target_unit_pci_target_sm_wr_progress
pci_target_unit_pci_target_sm_wr_to_fifo
pci_target_unit_pcit_if_pcir_fifo_control_in_637
pci_target_unit_pcit_if_pcir_fifo_data_in
pci_target_unit_pcit_if_pcir_fifo_data_in_766
pci_target_unit_pcit_if_pcir_fifo_data_in_767
pci_target_unit_pcit_if_pcir_fifo_data_in_768
pci_target_unit_pcit_if_pcir_fifo_data_in_769
pci_target_unit_pcit_if_pcir_fifo_data_in_770
pci_target_unit_pcit_if_pcir_fifo_data_in_771
pci_target_unit_pcit_if_pcir_fifo_data_in_772
pci_target_unit_pcit_if_pcir_fifo_data_in_773
pci_target_unit_pcit_if_pcir_fifo_data_in_774
pci_target_unit_pcit_if_pcir_fifo_data_in_775
pci_target_unit_pcit_if_pcir_fifo_data_in_776
pci_target_unit_pcit_if_pcir_fifo_data_in_777
pci_target_unit_pcit_if_pcir_fifo_data_in_778
pci_target_unit_pcit_if_pcir_fifo_data_in_779
pci_target_unit_pcit_if_pcir_fifo_data_in_780
pci_target_unit_pcit_if_pcir_fifo_data_in_781
pci_target_unit_pcit_if_pcir_fifo_data_in_782
pci_target_unit_pcit_if_pcir_fifo_data_in_783
pci_target_unit_pcit_if_pcir_fifo_data_in_784
pci_target_unit_pcit_if_pcir_fifo_data_in_785
pci_target_unit_pcit_if_pcir_fifo_data_in_786
pci_target_unit_pcit_if_pcir_fifo_data_in_787
pci_target_unit_pcit_if_pcir_fifo_data_in_788
pci_target_unit_pcit_if_pcir_fifo_data_in_789
pci_target_unit_pcit_if_pcir_fifo_data_in_790
pci_target_unit_pcit_if_pcir_fifo_data_in_791
pci_target_unit_pcit_if_pcir_fifo_data_in_792
pci_target_unit_pcit_if_pcir_fifo_data_in_793
pci_target_unit_pcit_if_pcir_fifo_data_in_794
pci_target_unit_pcit_if_pcir_fifo_data_in_795
pci_target_unit_pcit_if_pcir_fifo_data_in_796
pci_target_unit_pcit_if_req_req_pending_in
pci_target_unit_pcit_if_strd_addr_in_687
pci_target_unit_pcit_if_strd_addr_in_688
pci_target_unit_pcit_if_strd_addr_in_689
pci_target_unit_pcit_if_strd_addr_in_690
pci_target_unit_pcit_if_strd_addr_in_691
pci_target_unit_pcit_if_strd_addr_in_692
pci_target_unit_pcit_if_strd_addr_in_693
pci_target_unit_pcit_if_strd_addr_in_694
pci_target_unit_pcit_if_strd_addr_in_695
pci_target_unit_pcit_if_strd_addr_in_696
pci_target_unit_pcit_if_strd_addr_in_698
pci_target_unit_pcit_if_strd_addr_in_699
pci_target_unit_pcit_if_strd_addr_in_700
pci_target_unit_pcit_if_strd_addr_in_701
pci_target_unit_pcit_if_strd_addr_in_702
pci_target_unit_pcit_if_strd_addr_in_703
pci_target_unit_pcit_if_strd_addr_in_704
pci_target_unit_pcit_if_strd_addr_in_705
pci_target_unit_pcit_if_strd_addr_in_706
pci_target_unit_pcit_if_strd_addr_in_707
pci_target_unit_pcit_if_strd_addr_in_708
pci_target_unit_pcit_if_strd_addr_in_709
pci_target_unit_pcit_if_strd_addr_in_710
pci_target_unit_pcit_if_strd_addr_in_711
pci_target_unit_pcit_if_strd_addr_in_712
pci_target_unit_pcit_if_strd_addr_in_713
pci_target_unit_pcit_if_strd_addr_in_714
pci_target_unit_pcit_if_strd_addr_in_715
pci_target_unit_pcit_if_strd_addr_in_716
pci_target_unit_pcit_if_strd_bc_in
pci_target_unit_pcit_if_strd_bc_in_717
pci_target_unit_pcit_if_strd_bc_in_718
pci_target_unit_pcit_if_strd_bc_in_719
pci_target_unit_wbm_sm_pci_tar_burst_ok
pci_target_unit_wbm_sm_pci_tar_read_request
pci_target_unit_wbm_sm_pciw_fifo_addr_data_in
pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_50
pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_51
pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_52
pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_53
pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_54
pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_55
pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_56
pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_57
pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_58
pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_59
pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_60
pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_61
pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_62
pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_63
pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_64
pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_65
pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_66
pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_67
pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_68
pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_69
pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_70
pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_71
pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_72
pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_73
pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_74
pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_75
pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_76
pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_77
pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_78
pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_79
pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_80
pci_target_unit_wbm_sm_pciw_fifo_cbe_in
pci_target_unit_wbm_sm_pciw_fifo_cbe_in_81
pci_target_unit_wbm_sm_pciw_fifo_cbe_in_82
pci_target_unit_wbm_sm_pciw_fifo_cbe_in_83
pci_target_unit_wbm_sm_pciw_fifo_control_in
pci_target_unit_wbm_sm_pciw_fifo_control_in_84
pci_target_unit_wbm_sm_pciw_fifo_control_in_85
pci_target_unit_wbm_sm_pciw_fifo_control_in_86
pci_target_unit_wishbone_master_addr_into_cnt_reg
pci_target_unit_wishbone_master_bc_register_reg_0__Q
pci_target_unit_wishbone_master_bc_register_reg_1__Q
pci_target_unit_wishbone_master_bc_register_reg_2__Q
pci_target_unit_wishbone_master_bc_register_reg_3__Q
pci_target_unit_wishbone_master_burst_chopped
pci_target_unit_wishbone_master_burst_chopped_delayed
pci_target_unit_wishbone_master_burst_chopped_delayed_reg_Q
pci_target_unit_wishbone_master_c_state_0_
pci_target_unit_wishbone_master_c_state_1_
pci_target_unit_wishbone_master_c_state_2_
pci_target_unit_wishbone_master_first_data_is_burst_reg
pci_target_unit_wishbone_master_first_wb_data_access
pci_target_unit_wishbone_master_read_bound
pci_target_unit_wishbone_master_read_count_0_
pci_target_unit_wishbone_master_read_count_1_
pci_target_unit_wishbone_master_read_count_reg_2__Q
pci_target_unit_wishbone_master_reset_rty_cnt
pci_target_unit_wishbone_master_reset_rty_cnt_reg_Q
pci_target_unit_wishbone_master_retried
pci_target_unit_wishbone_master_rty_counter_0_
pci_target_unit_wishbone_master_rty_counter_1_
pci_target_unit_wishbone_master_rty_counter_3_
pci_target_unit_wishbone_master_rty_counter_4_
pci_target_unit_wishbone_master_rty_counter_5_
pci_target_unit_wishbone_master_rty_counter_6_
pci_target_unit_wishbone_master_rty_counter_7_
pci_target_unit_wishbone_master_wb_cyc_o_reg_Q
pciu_am1_in
pciu_am1_in_518
pciu_am1_in_521
pciu_am1_in_522
pciu_am1_in_523
pciu_am1_in_524
pciu_am1_in_525
pciu_am1_in_526
pciu_am1_in_527
pciu_am1_in_528
pciu_am1_in_529
pciu_am1_in_530
pciu_am1_in_531
pciu_am1_in_533
pciu_am1_in_536
pciu_am1_in_537
pciu_am1_in_538
pciu_am1_in_539
pciu_am1_in_540
pciu_bar0_in
pciu_bar0_in_361
pciu_bar0_in_362
pciu_bar0_in_363
pciu_bar0_in_364
pciu_bar0_in_365
pciu_bar0_in_366
pciu_bar0_in_367
pciu_bar0_in_368
pciu_bar0_in_369
pciu_bar0_in_372
pciu_bar0_in_373
pciu_bar0_in_374
pciu_bar0_in_375
pciu_bar0_in_376
pciu_bar0_in_377
pciu_bar0_in_378
pciu_bar0_in_379
pciu_bar1_in_380
pciu_bar1_in_382
pciu_bar1_in_383
pciu_bar1_in_384
pciu_bar1_in_385
pciu_bar1_in_386
pciu_bar1_in_388
pciu_bar1_in_389
pciu_bar1_in_390
pciu_bar1_in_391
pciu_bar1_in_392
pciu_bar1_in_395
pciu_bar1_in_396
pciu_bar1_in_398
pciu_bar1_in_399
pciu_bar1_in_400
pciu_bar1_in_401
pciu_bar1_in_402
pciu_cache_lsize_not_zero_in
pciu_pciif_bckp_stop_in
pciu_pciif_idsel_reg_in
pciu_pref_en_in_320
wbm_cyc_o_1378
wbs_ack_o_1307
wbs_err_o_1309
wbs_wbb3_2_wbb2_dat_o_i
wbs_wbb3_2_wbb2_dat_o_i_100
wbs_wbb3_2_wbb2_dat_o_i_101
wbs_wbb3_2_wbb2_dat_o_i_103
wbs_wbb3_2_wbb2_dat_o_i_104
wbs_wbb3_2_wbb2_dat_o_i_105
wbs_wbb3_2_wbb2_dat_o_i_106
wbs_wbb3_2_wbb2_dat_o_i_107
wbs_wbb3_2_wbb2_dat_o_i_108
wbs_wbb3_2_wbb2_dat_o_i_109
wbs_wbb3_2_wbb2_dat_o_i_110
wbs_wbb3_2_wbb2_dat_o_i_111
wbs_wbb3_2_wbb2_dat_o_i_112
wbs_wbb3_2_wbb2_dat_o_i_113
wbs_wbb3_2_wbb2_dat_o_i_114
wbs_wbb3_2_wbb2_dat_o_i_115
wbs_wbb3_2_wbb2_dat_o_i_116
wbs_wbb3_2_wbb2_dat_o_i_117
wbs_wbb3_2_wbb2_dat_o_i_118
wbs_wbb3_2_wbb2_dat_o_i_119
wbs_wbb3_2_wbb2_dat_o_i_120
wbs_wbb3_2_wbb2_dat_o_i_121
wbs_wbb3_2_wbb2_dat_o_i_122
wbs_wbb3_2_wbb2_dat_o_i_123
wbs_wbb3_2_wbb2_dat_o_i_124
wbs_wbb3_2_wbb2_dat_o_i_125
wbs_wbb3_2_wbb2_dat_o_i_126
wbs_wbb3_2_wbb2_dat_o_i_127
wbs_wbb3_2_wbb2_dat_o_i_128
wbs_wbb3_2_wbb2_dat_o_i_129
wbs_wbb3_2_wbb2_dat_o_i_130
wbu_addr_in
wbu_addr_in_250
wbu_addr_in_251
wbu_addr_in_252
wbu_addr_in_253
wbu_addr_in_254
wbu_addr_in_255
wbu_addr_in_256
wbu_addr_in_257
wbu_addr_in_258
wbu_addr_in_259
wbu_addr_in_260
wbu_addr_in_261
wbu_addr_in_262
wbu_addr_in_263
wbu_addr_in_264
wbu_addr_in_265
wbu_addr_in_266
wbu_addr_in_267
wbu_addr_in_268
wbu_addr_in_269
wbu_addr_in_270
wbu_addr_in_271
wbu_addr_in_272
wbu_addr_in_273
wbu_addr_in_274
wbu_addr_in_275
wbu_addr_in_276
wbu_addr_in_277
wbu_addr_in_278
wbu_addr_in_279
wbu_addr_in_280
wbu_am1_in
wbu_am2_in
wbu_bar1_in
wbu_bar2_in
wbu_cache_line_size_in_206
wbu_cache_line_size_in_207
wbu_cache_line_size_in_208
wbu_cache_line_size_in_209
wbu_cache_line_size_in_210
wbu_cache_line_size_in_211
wbu_latency_tim_val_in_247
wbu_map_in_131
wbu_map_in_132
wbu_mrl_en_in_141
wbu_mrl_en_in_142
wbu_pci_drcomp_pending_in
wbu_pciif_devsel_reg_in
wbu_pref_en_in_136
wbu_pref_en_in_137
wbu_sel_in_312
wbu_sel_in_313
wbu_sel_in_314
wbu_wb_init_complete_in
wishbone_slave_unit_del_sync_addr_out_reg_0__Q
wishbone_slave_unit_del_sync_addr_out_reg_10__Q
wishbone_slave_unit_del_sync_addr_out_reg_11__Q
wishbone_slave_unit_del_sync_addr_out_reg_12__Q
wishbone_slave_unit_del_sync_addr_out_reg_13__Q
wishbone_slave_unit_del_sync_addr_out_reg_14__Q
wishbone_slave_unit_del_sync_addr_out_reg_15__Q
wishbone_slave_unit_del_sync_addr_out_reg_16__Q
wishbone_slave_unit_del_sync_addr_out_reg_17__Q
wishbone_slave_unit_del_sync_addr_out_reg_18__Q
wishbone_slave_unit_del_sync_addr_out_reg_19__Q
wishbone_slave_unit_del_sync_addr_out_reg_1__Q
wishbone_slave_unit_del_sync_addr_out_reg_20__Q
wishbone_slave_unit_del_sync_addr_out_reg_21__Q
wishbone_slave_unit_del_sync_addr_out_reg_22__Q
wishbone_slave_unit_del_sync_addr_out_reg_23__Q
wishbone_slave_unit_del_sync_addr_out_reg_24__Q
wishbone_slave_unit_del_sync_addr_out_reg_25__Q
wishbone_slave_unit_del_sync_addr_out_reg_26__Q
wishbone_slave_unit_del_sync_addr_out_reg_27__Q
wishbone_slave_unit_del_sync_addr_out_reg_28__Q
wishbone_slave_unit_del_sync_addr_out_reg_29__Q
wishbone_slave_unit_del_sync_addr_out_reg_2__Q
wishbone_slave_unit_del_sync_addr_out_reg_30__Q
wishbone_slave_unit_del_sync_addr_out_reg_31__Q
wishbone_slave_unit_del_sync_addr_out_reg_3__Q
wishbone_slave_unit_del_sync_addr_out_reg_4__Q
wishbone_slave_unit_del_sync_addr_out_reg_5__Q
wishbone_slave_unit_del_sync_addr_out_reg_6__Q
wishbone_slave_unit_del_sync_addr_out_reg_7__Q
wishbone_slave_unit_del_sync_addr_out_reg_8__Q
wishbone_slave_unit_del_sync_addr_out_reg_9__Q
wishbone_slave_unit_del_sync_comp_comp_pending_reg_Q
wishbone_slave_unit_del_sync_comp_cycle_count_0_
wishbone_slave_unit_del_sync_comp_cycle_count_10_
wishbone_slave_unit_del_sync_comp_cycle_count_1_
wishbone_slave_unit_del_sync_comp_cycle_count_2_
wishbone_slave_unit_del_sync_comp_cycle_count_3_
wishbone_slave_unit_del_sync_comp_cycle_count_4_
wishbone_slave_unit_del_sync_comp_cycle_count_5_
wishbone_slave_unit_del_sync_comp_cycle_count_6_
wishbone_slave_unit_del_sync_comp_cycle_count_7_
wishbone_slave_unit_del_sync_comp_cycle_count_reg_16__Q
wishbone_slave_unit_del_sync_comp_done_reg_clr
wishbone_slave_unit_del_sync_comp_done_reg_clr_reg_Q
wishbone_slave_unit_del_sync_comp_done_reg_main
wishbone_slave_unit_del_sync_comp_flush_out
wishbone_slave_unit_del_sync_comp_req_pending_reg_Q
wishbone_slave_unit_del_sync_comp_rty_exp_reg
wishbone_slave_unit_del_sync_req_comp_pending
wishbone_slave_unit_del_sync_req_comp_pending_sample
wishbone_slave_unit_del_sync_req_comp_pending_sample_reg_Q
wishbone_slave_unit_del_sync_req_done_reg
wishbone_slave_unit_del_sync_req_done_reg_reg_Q
wishbone_slave_unit_del_sync_req_rty_exp_clr
wishbone_slave_unit_del_sync_req_rty_exp_reg
wishbone_slave_unit_del_sync_sync_comp_done
wishbone_slave_unit_del_sync_sync_comp_req_pending
wishbone_slave_unit_del_sync_sync_req_comp_pending
wishbone_slave_unit_del_sync_sync_req_rty_exp
wishbone_slave_unit_del_sync_we_out_reg_Q
wishbone_slave_unit_delayed_write_data_comp_wdata_out_100
wishbone_slave_unit_delayed_write_data_comp_wdata_out_101
wishbone_slave_unit_delayed_write_data_comp_wdata_out_70
wishbone_slave_unit_delayed_write_data_comp_wdata_out_71
wishbone_slave_unit_delayed_write_data_comp_wdata_out_73
wishbone_slave_unit_delayed_write_data_comp_wdata_out_75
wishbone_slave_unit_delayed_write_data_comp_wdata_out_76
wishbone_slave_unit_delayed_write_data_comp_wdata_out_80
wishbone_slave_unit_delayed_write_data_comp_wdata_out_81
wishbone_slave_unit_delayed_write_data_comp_wdata_out_83
wishbone_slave_unit_delayed_write_data_comp_wdata_out_84
wishbone_slave_unit_delayed_write_data_comp_wdata_out_85
wishbone_slave_unit_delayed_write_data_comp_wdata_out_86
wishbone_slave_unit_delayed_write_data_comp_wdata_out_87
wishbone_slave_unit_delayed_write_data_comp_wdata_out_88
wishbone_slave_unit_delayed_write_data_comp_wdata_out_90
wishbone_slave_unit_delayed_write_data_comp_wdata_out_91
wishbone_slave_unit_delayed_write_data_comp_wdata_out_93
wishbone_slave_unit_delayed_write_data_comp_wdata_out_96
wishbone_slave_unit_delayed_write_data_comp_wdata_out_97
wishbone_slave_unit_delayed_write_data_comp_wdata_out_98
wishbone_slave_unit_delayed_write_data_comp_wdata_out_99
wishbone_slave_unit_fifos_inGreyCount_0_
wishbone_slave_unit_fifos_inGreyCount_reg_0__Q
wishbone_slave_unit_fifos_inGreyCount_reg_1__Q
wishbone_slave_unit_fifos_inGreyCount_reg_2__Q
wishbone_slave_unit_fifos_outGreyCount_0_
wishbone_slave_unit_fifos_outGreyCount_1_
wishbone_slave_unit_fifos_outGreyCount_2_
wishbone_slave_unit_fifos_pci_clk_inGreyCount_0_
wishbone_slave_unit_fifos_pci_clk_inGreyCount_1_
wishbone_slave_unit_fifos_pci_clk_inGreyCount_2_
wishbone_slave_unit_fifos_pci_clk_inGreyCount_reg_2__Q
wishbone_slave_unit_fifos_pci_clk_sync_inGreyCount
wishbone_slave_unit_fifos_pci_clk_sync_inGreyCount_49
wishbone_slave_unit_fifos_pci_clk_sync_inGreyCount_50
wishbone_slave_unit_fifos_wbr_be_in_264
wishbone_slave_unit_fifos_wbr_be_in_265
wishbone_slave_unit_fifos_wbr_be_in_266
wishbone_slave_unit_fifos_wbr_control_in
wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_0_
wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_1_
wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_2_
wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_0_
wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_1_
wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_2_
wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_3_
wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg_0__Q
wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg_1__Q
wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg_2__Q
wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg_3__Q
wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg_0__Q
wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg_1__Q
wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg_2__Q
wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg_3__Q
wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_sync_wgrey_addr
wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_sync_wgrey_addr_45
wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_sync_wgrey_addr_46
wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_sync_wgrey_addr_47
wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_0_
wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_1_
wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_2_
wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_3_
wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg_0__Q
wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg_1__Q
wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg_2__Q
wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg_3__Q
wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_0_
wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_1_
wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_2_
wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_3_
wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_0_
wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg_0__Q
wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg_1__Q
wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg_2__Q
wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg_3__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__43
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__46
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__47
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__51
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__59
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__62
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__67
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_11__466
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_12__484
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_13__509
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_13__522
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_13__531
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_13__532
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_13__536
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_13__544
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_15__622
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_3__177
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_3__178
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_3__183
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__258
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__271
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_8__330
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_8__342
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__358
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__360
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__374
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__376
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__377
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__380
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__0__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__12__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__14__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__18__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__20__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__21__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__22__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__23__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__24__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__25__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__26__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__28__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__29__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__37__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__4__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__6__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__7__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__8__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__9__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__10__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__11__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__12__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__15__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__16__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__18__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__19__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__21__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__22__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__23__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__25__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__26__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__28__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__29__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__2__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__30__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__37__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__3__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__4__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__5__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__7__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__8__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__0__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__12__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__15__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__18__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__1__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__21__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__22__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__23__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__24__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__25__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__27__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__28__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__29__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__2__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__31__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__36__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__37__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__3__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__4__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__5__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__6__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__8__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__9__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__10__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__11__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__12__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__17__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__18__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__1__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__20__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__21__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__24__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__27__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__29__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__31__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__37__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__3__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__4__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__5__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__7__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__8__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__9__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__10__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__12__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__14__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__15__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__18__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__19__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__1__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__20__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__21__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__22__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__23__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__24__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__25__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__26__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__28__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__29__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__2__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__30__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__37__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__5__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__6__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__8__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__10__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__11__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__12__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__14__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__17__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__19__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__1__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__20__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__21__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__23__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__25__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__27__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__28__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__29__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__3__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__7__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__9__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__10__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__12__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__14__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__15__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__18__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__19__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__1__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__20__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__22__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__23__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__24__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__25__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__27__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__29__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__30__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__37__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__5__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__6__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__7__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__8__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__11__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__12__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__15__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__16__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__18__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__20__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__21__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__22__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__24__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__26__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__27__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__28__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__29__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__2__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__30__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__37__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__5__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__6__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__8__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__11__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__12__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__15__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__16__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__17__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__1__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__20__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__21__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__22__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__23__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__24__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__26__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__27__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__29__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__30__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__36__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__37__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__3__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__4__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__5__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__6__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__7__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__9__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__0__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__12__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__13__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__15__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__16__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__17__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__1__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__21__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__23__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__24__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__25__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__27__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__28__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__29__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__2__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__31__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__3__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__4__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__7__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__9__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__10__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__12__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__16__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__17__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__18__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__1__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__20__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__21__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__23__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__24__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__25__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__26__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__27__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__28__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__29__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__30__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__37__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__3__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__4__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__5__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__7__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__8__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__0__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__11__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__12__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__13__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__15__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__16__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__17__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__19__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__1__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__21__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__22__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__23__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__24__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__25__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__27__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__28__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__29__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__30__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__31__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__37__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__3__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__6__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__7__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__8__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__9__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__10__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__12__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__16__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__17__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__18__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__19__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__1__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__23__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__24__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__25__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__27__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__28__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__29__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__30__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__37__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__6__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__7__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__8__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__10__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__11__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__12__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__16__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__17__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__19__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__21__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__23__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__25__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__28__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__29__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__3__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__5__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__6__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__8__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__12__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__16__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__18__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__19__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__1__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__20__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__21__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__22__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__23__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__24__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__25__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__27__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__28__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__29__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__2__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__30__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__31__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__37__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__3__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__4__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__5__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__6__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__8__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__9__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__10__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__11__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__14__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__15__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__16__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__17__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__18__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__19__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__21__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__23__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__25__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__26__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__27__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__29__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__2__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__30__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__37__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__3__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__5__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__7__Q
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__9__Q
wishbone_slave_unit_fifos_wbr_whole_waddr
wishbone_slave_unit_fifos_wbr_whole_waddr_104
wishbone_slave_unit_fifos_wbr_whole_waddr_105
wishbone_slave_unit_fifos_wbr_whole_waddr_106
wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_0_
wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_1_
wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_2_
wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_3_
wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_0_
wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_1_
wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_2_
wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_3_
wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_sync_wgrey_next
wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_sync_wgrey_next_70
wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_sync_wgrey_next_71
wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_sync_wgrey_next_72
wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_0_
wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_1_
wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_2_
wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_3_
wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_addr_reg_0__Q
wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_addr_reg_1__Q
wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_addr_reg_2__Q
wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_addr_reg_3__Q
wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_minus1_reg_0__Q
wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_minus1_reg_1__Q
wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_minus1_reg_2__Q
wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_minus1_reg_3__Q
wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_0_
wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_1_
wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_2_
wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_3_
wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_0_
wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_1_
wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_2_
wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_3_
wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_sync_rgrey_minus1
wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_sync_rgrey_minus_93
wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_sync_rgrey_minus_94
wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_sync_rgrey_minus_95
wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_0_
wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_1_
wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_2_
wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_3_
wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_0_
wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_1_
wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_2_
wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_3_
wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_33__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_14__582
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_15__621
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_7__309
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__0__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__10__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__11__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__12__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__13__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__14__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__15__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__16__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__17__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__19__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__1__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__20__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__21__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__22__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__23__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__24__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__25__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__26__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__27__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__28__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__29__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__2__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__31__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__32__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__33__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__34__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__35__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__3__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__5__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__6__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__8__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__9__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__0__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__10__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__11__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__13__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__14__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__15__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__16__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__17__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__19__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__1__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__20__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__21__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__22__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__23__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__24__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__26__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__27__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__28__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__29__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__2__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__30__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__31__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__32__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__33__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__34__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__35__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__5__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__6__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__9__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__0__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__10__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__11__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__12__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__13__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__14__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__15__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__16__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__17__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__18__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__19__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__1__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__20__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__22__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__23__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__24__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__25__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__26__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__27__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__28__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__29__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__31__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__33__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__3__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__5__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__6__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__7__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__8__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__9__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__0__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__10__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__11__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__12__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__13__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__14__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__15__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__16__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__17__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__18__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__19__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__20__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__21__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__22__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__23__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__24__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__25__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__26__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__27__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__28__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__29__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__2__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__30__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__31__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__33__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__34__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__4__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__5__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__6__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__8__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__9__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__0__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__12__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__13__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__14__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__15__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__16__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__17__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__18__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__19__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__1__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__20__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__21__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__23__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__24__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__25__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__26__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__27__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__28__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__29__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__30__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__31__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__32__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__33__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__34__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__35__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__3__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__4__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__5__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__6__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__8__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__0__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__10__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__11__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__12__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__13__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__14__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__15__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__16__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__17__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__18__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__19__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__1__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__20__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__21__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__22__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__23__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__24__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__25__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__26__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__27__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__28__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__29__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__2__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__30__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__31__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__33__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__34__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__35__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__36__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__4__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__5__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__6__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__7__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__8__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__9__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__0__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__10__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__12__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__13__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__14__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__15__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__16__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__17__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__18__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__19__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__1__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__20__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__21__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__23__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__24__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__26__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__27__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__28__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__29__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__30__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__31__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__32__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__33__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__34__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__35__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__36__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__3__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__4__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__5__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__6__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__10__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__11__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__12__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__13__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__14__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__15__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__16__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__17__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__19__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__20__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__21__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__22__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__23__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__24__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__25__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__26__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__27__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__28__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__2__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__31__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__33__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__3__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__5__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__6__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__7__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__8__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__9__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__10__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__11__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__12__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__13__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__14__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__15__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__16__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__17__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__19__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__20__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__21__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__22__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__23__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__24__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__25__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__26__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__27__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__28__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__29__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__2__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__30__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__31__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__33__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__36__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__3__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__5__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__6__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__7__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__8__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__9__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__10__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__12__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__13__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__14__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__15__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__16__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__17__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__19__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__20__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__22__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__23__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__24__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__25__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__26__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__27__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__28__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__29__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__2__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__30__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__31__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__33__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__34__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__36__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__3__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__4__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__5__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__6__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__7__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__8__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__0__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__10__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__11__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__13__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__14__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__15__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__16__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__17__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__19__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__1__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__20__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__21__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__22__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__23__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__24__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__26__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__27__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__28__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__29__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__2__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__31__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__32__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__33__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__35__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__5__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__6__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__8__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__9__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__10__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__12__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__13__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__14__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__15__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__16__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__17__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__19__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__20__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__21__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__23__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__24__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__25__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__26__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__27__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__28__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__29__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__30__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__31__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__33__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__34__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__35__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__3__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__4__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__5__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__6__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__7__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__8__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__0__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__11__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__14__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__16__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__17__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__19__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__1__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__20__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__21__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__22__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__23__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__24__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__26__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__27__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__28__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__29__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__2__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__30__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__32__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__33__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__35__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__3__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__4__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__5__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__6__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__9__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__0__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__10__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__11__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__14__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__16__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__17__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__18__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__19__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__1__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__20__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__21__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__22__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__23__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__24__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__27__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__28__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__2__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__30__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__32__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__33__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__35__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__36__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__3__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__5__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__6__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__9__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__0__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__10__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__11__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__12__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__13__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__14__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__15__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__16__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__17__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__18__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__19__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__1__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__20__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__22__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__23__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__24__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__25__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__26__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__27__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__28__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__29__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__30__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__31__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__33__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__36__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__3__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__5__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__6__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__7__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__8__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__9__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__0__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__10__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__11__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__13__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__14__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__15__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__16__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__17__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__18__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__19__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__1__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__20__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__21__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__22__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__23__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__24__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__26__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__27__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__28__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__29__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__2__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__30__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__31__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__32__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__33__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__34__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__35__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__3__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__5__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__6__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__7__Q
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__9__Q
wishbone_slave_unit_fifos_wbw_inTransactionCount_0_
wishbone_slave_unit_fifos_wbw_inTransactionCount_1_
wishbone_slave_unit_fifos_wbw_inTransactionCount_reg_0__Q
wishbone_slave_unit_fifos_wbw_inTransactionCount_reg_1__Q
wishbone_slave_unit_fifos_wbw_inTransactionCount_reg_2__Q
wishbone_slave_unit_fifos_wbw_outTransactionCount_0_
wishbone_slave_unit_fifos_wbw_outTransactionCount_1_
wishbone_slave_unit_fifos_wbw_outTransactionCount_reg_0__Q
wishbone_slave_unit_fifos_wbw_outTransactionCount_reg_1__Q
wishbone_slave_unit_fifos_wbw_outTransactionCount_reg_2__Q
wishbone_slave_unit_fifos_wbw_whole_waddr
wishbone_slave_unit_fifos_wbw_whole_waddr_55
wishbone_slave_unit_fifos_wbw_whole_waddr_56
wishbone_slave_unit_fifos_wbw_whole_waddr_57
wishbone_slave_unit_pci_initiator_if_current_byte_address
wishbone_slave_unit_pci_initiator_if_current_byte_address_36
wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_29__Q
wishbone_slave_unit_pci_initiator_if_data_source
wishbone_slave_unit_pci_initiator_if_del_read_req
wishbone_slave_unit_pci_initiator_if_del_write_req
wishbone_slave_unit_pci_initiator_if_err_recovery
wishbone_slave_unit_pci_initiator_if_intermediate_be_reg_2__Q
wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_0__Q
wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_10__Q
wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_11__Q
wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_13__Q
wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_14__Q
wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_15__Q
wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_16__Q
wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_17__Q
wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_18__Q
wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_19__Q
wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_1__Q
wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_20__Q
wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_21__Q
wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_23__Q
wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_24__Q
wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_25__Q
wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_27__Q
wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_28__Q
wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_29__Q
wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_30__Q
wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_31__Q
wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_3__Q
wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_4__Q
wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_5__Q
wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_6__Q
wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_7__Q
wishbone_slave_unit_pci_initiator_if_read_count_0_
wishbone_slave_unit_pci_initiator_if_tabort_received_out_reg_Q
wishbone_slave_unit_pci_initiator_sm_cur_state_0_
wishbone_slave_unit_pci_initiator_sm_cur_state_1_
wishbone_slave_unit_pci_initiator_sm_cur_state_2_
wishbone_slave_unit_pci_initiator_sm_cur_state_3_
wishbone_slave_unit_pci_initiator_sm_decode_count_0_
wishbone_slave_unit_pci_initiator_sm_decode_count_1_
wishbone_slave_unit_pci_initiator_sm_decode_count_2_
wishbone_slave_unit_pci_initiator_sm_latency_timer_4_
wishbone_slave_unit_pci_initiator_sm_latency_timer_5_
wishbone_slave_unit_pci_initiator_sm_mabort1
wishbone_slave_unit_pci_initiator_sm_rdata_selector
wishbone_slave_unit_pci_initiator_sm_rdata_selector_14
wishbone_slave_unit_pcim_if_del_burst_in
wishbone_slave_unit_pcim_if_del_req_in
wishbone_slave_unit_pcim_if_del_we_in
wishbone_slave_unit_pcim_if_wbw_addr_data_in
wishbone_slave_unit_pcim_if_wbw_addr_data_in_384
wishbone_slave_unit_pcim_if_wbw_addr_data_in_385
wishbone_slave_unit_pcim_if_wbw_addr_data_in_386
wishbone_slave_unit_pcim_if_wbw_addr_data_in_387
wishbone_slave_unit_pcim_if_wbw_addr_data_in_388
wishbone_slave_unit_pcim_if_wbw_addr_data_in_389
wishbone_slave_unit_pcim_if_wbw_addr_data_in_390
wishbone_slave_unit_pcim_if_wbw_addr_data_in_391
wishbone_slave_unit_pcim_if_wbw_addr_data_in_392
wishbone_slave_unit_pcim_if_wbw_addr_data_in_393
wishbone_slave_unit_pcim_if_wbw_addr_data_in_394
wishbone_slave_unit_pcim_if_wbw_addr_data_in_395
wishbone_slave_unit_pcim_if_wbw_addr_data_in_396
wishbone_slave_unit_pcim_if_wbw_addr_data_in_397
wishbone_slave_unit_pcim_if_wbw_addr_data_in_398
wishbone_slave_unit_pcim_if_wbw_addr_data_in_399
wishbone_slave_unit_pcim_if_wbw_addr_data_in_400
wishbone_slave_unit_pcim_if_wbw_addr_data_in_401
wishbone_slave_unit_pcim_if_wbw_addr_data_in_402
wishbone_slave_unit_pcim_if_wbw_addr_data_in_403
wishbone_slave_unit_pcim_if_wbw_addr_data_in_404
wishbone_slave_unit_pcim_if_wbw_addr_data_in_405
wishbone_slave_unit_pcim_if_wbw_addr_data_in_406
wishbone_slave_unit_pcim_if_wbw_addr_data_in_407
wishbone_slave_unit_pcim_if_wbw_addr_data_in_408
wishbone_slave_unit_pcim_if_wbw_addr_data_in_409
wishbone_slave_unit_pcim_if_wbw_addr_data_in_410
wishbone_slave_unit_pcim_if_wbw_addr_data_in_411
wishbone_slave_unit_pcim_if_wbw_addr_data_in_412
wishbone_slave_unit_pcim_if_wbw_addr_data_in_413
wishbone_slave_unit_pcim_if_wbw_addr_data_in_414
wishbone_slave_unit_pcim_if_wbw_cbe_in_416
wishbone_slave_unit_pcim_sm_be_in_557
wishbone_slave_unit_pcim_sm_be_in_558
wishbone_slave_unit_pcim_sm_be_in_559
wishbone_slave_unit_pcim_sm_data_in
wishbone_slave_unit_pcim_sm_data_in_635
wishbone_slave_unit_pcim_sm_data_in_636
wishbone_slave_unit_pcim_sm_data_in_637
wishbone_slave_unit_pcim_sm_data_in_638
wishbone_slave_unit_pcim_sm_data_in_639
wishbone_slave_unit_pcim_sm_data_in_640
wishbone_slave_unit_pcim_sm_data_in_641
wishbone_slave_unit_pcim_sm_data_in_643
wishbone_slave_unit_pcim_sm_data_in_644
wishbone_slave_unit_pcim_sm_data_in_645
wishbone_slave_unit_pcim_sm_data_in_646
wishbone_slave_unit_pcim_sm_data_in_647
wishbone_slave_unit_pcim_sm_data_in_648
wishbone_slave_unit_pcim_sm_data_in_649
wishbone_slave_unit_pcim_sm_data_in_650
wishbone_slave_unit_pcim_sm_data_in_651
wishbone_slave_unit_pcim_sm_data_in_652
wishbone_slave_unit_pcim_sm_data_in_653
wishbone_slave_unit_pcim_sm_data_in_654
wishbone_slave_unit_pcim_sm_data_in_655
wishbone_slave_unit_pcim_sm_data_in_657
wishbone_slave_unit_pcim_sm_data_in_658
wishbone_slave_unit_pcim_sm_data_in_659
wishbone_slave_unit_pcim_sm_data_in_660
wishbone_slave_unit_pcim_sm_data_in_661
wishbone_slave_unit_pcim_sm_data_in_662
wishbone_slave_unit_pcim_sm_data_in_663
wishbone_slave_unit_pcim_sm_data_in_664
wishbone_slave_unit_pcim_sm_data_in_665
wishbone_slave_unit_pcim_sm_rdy_in
wishbone_slave_unit_wbs_sm_del_req_pending_in
wishbone_slave_unit_wbs_sm_wbr_control_in
wishbone_slave_unit_wbs_sm_wbr_control_in_190
wishbone_slave_unit_wishbone_slave_async_reset_as_wbr_flush_async_reset_data_out_reg_Q
wishbone_slave_unit_wishbone_slave_c_state
wishbone_slave_unit_wishbone_slave_c_state_1
wishbone_slave_unit_wishbone_slave_c_state_2
wishbone_slave_unit_wishbone_slave_d_incoming_reg_0__Q
wishbone_slave_unit_wishbone_slave_d_incoming_reg_10__Q
wishbone_slave_unit_wishbone_slave_d_incoming_reg_11__Q
wishbone_slave_unit_wishbone_slave_d_incoming_reg_12__Q
wishbone_slave_unit_wishbone_slave_d_incoming_reg_13__Q
wishbone_slave_unit_wishbone_slave_d_incoming_reg_14__Q
wishbone_slave_unit_wishbone_slave_d_incoming_reg_15__Q
wishbone_slave_unit_wishbone_slave_d_incoming_reg_16__Q
wishbone_slave_unit_wishbone_slave_d_incoming_reg_17__Q
wishbone_slave_unit_wishbone_slave_d_incoming_reg_18__Q
wishbone_slave_unit_wishbone_slave_d_incoming_reg_19__Q
wishbone_slave_unit_wishbone_slave_d_incoming_reg_1__Q
wishbone_slave_unit_wishbone_slave_d_incoming_reg_20__Q
wishbone_slave_unit_wishbone_slave_d_incoming_reg_21__Q
wishbone_slave_unit_wishbone_slave_d_incoming_reg_22__Q
wishbone_slave_unit_wishbone_slave_d_incoming_reg_23__Q
wishbone_slave_unit_wishbone_slave_d_incoming_reg_24__Q
wishbone_slave_unit_wishbone_slave_d_incoming_reg_25__Q
wishbone_slave_unit_wishbone_slave_d_incoming_reg_26__Q
wishbone_slave_unit_wishbone_slave_d_incoming_reg_27__Q
wishbone_slave_unit_wishbone_slave_d_incoming_reg_28__Q
wishbone_slave_unit_wishbone_slave_d_incoming_reg_29__Q
wishbone_slave_unit_wishbone_slave_d_incoming_reg_2__Q
wishbone_slave_unit_wishbone_slave_d_incoming_reg_30__Q
wishbone_slave_unit_wishbone_slave_d_incoming_reg_31__Q
wishbone_slave_unit_wishbone_slave_d_incoming_reg_3__Q
wishbone_slave_unit_wishbone_slave_d_incoming_reg_4__Q
wishbone_slave_unit_wishbone_slave_d_incoming_reg_6__Q
wishbone_slave_unit_wishbone_slave_d_incoming_reg_7__Q
wishbone_slave_unit_wishbone_slave_d_incoming_reg_8__Q
wishbone_slave_unit_wishbone_slave_d_incoming_reg_9__Q
wishbone_slave_unit_wishbone_slave_del_addr_hit
wishbone_slave_unit_wishbone_slave_del_completion_allow
wishbone_slave_unit_wishbone_slave_do_del_request
wishbone_slave_unit_wishbone_slave_img_hit_0_
wishbone_slave_unit_wishbone_slave_img_hit_1_
wishbone_slave_unit_wishbone_slave_img_hit_2_
wishbone_slave_unit_wishbone_slave_img_hit_3_
wishbone_slave_unit_wishbone_slave_img_hit_4_
wishbone_slave_unit_wishbone_slave_img_wallow
wishbone_slave_unit_wishbone_slave_wb_conf_hit
ec0/g65065_db
ec0/n_6289
ec0/g62632_db
ec0/g65092_db
ec0/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__27__Q
ec0/n_4299
ec0/n_6754
ec0/n_11814
ec0/g62936_sb
ec0/g64929_da
ec0/g64929_sb
ec0/n_12296
ec0/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__22__Q
ec0/n_3679
ec0/g62633_db
ec0/n_12075
ec0/g64994_sb
ec0/FE_OFN1144_n_6391
ec0/n_11937
ec0/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__5__Q
ec0/n_6430
ec0/g62564_db
ec0/n_13117
ec0/g62541_sb
ec0/g64944_sb
ec0/FE_OCPN1882_FE_OFN1454_n_12028
ec0/FE_OCP_RBN2083_n_10244
ec0/g62387_sb
ec0/n_12259
ec0/n_12689
ec0/n_12260
ec0/g65009_sb
ec0/g62966_sb
ec0/g62966_da
ec0/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__2__Q
ec0/n_4661
ec0/n_1688
ec0/g64022_p
ec0/n_1015
ec0/g65522_p2
ec0/wishbone_slave_unit_pci_initiator_sm_latency_timer_2_
ec0/n_4824
ec0/n_3045
ec0/n_3444
ec0/n_6987
ec0/FE_OFN1098_n_5592
ec0/g62123_db
ec0/n_5608
ec0/g62096_db
ec0/FE_OFN1096_n_5592
ec0/n_5607
ec0/g62097_db
ec0/n_5572
ec0/g62124_db
ec0/g62079_da
ec0/n_5617
ec0/g62090_db
ec0/n_5591
ec0/g62108_da
ec0/g62108_db
ec0/g62108_sb
ec0/n_2853
ec0/FE_OCPN1968_n_15445
ec0/FE_OFN1102_n_5592
ec0/configuration_wb_err_data_575
ec0/conf_wb_err_bc_in_847
ec0/n_1588
ec0/n_545
ec0/g61843_db
ec0/n_14390
ec0/n_13752
ec0/g61843_sb
ec0/n_13554
ec0/g53943_da
ec0/n_13502
ec0/g53943_db
ec0/n_13226
ec0/g59796_sb
ec0/g59796_db
ec0/g63533_sb
ec0/n_13224
ec0/g59799_sb
ec0/g54169_db
ec0/n_398
ec0/g54166_db
ec0/n_8673
ec0/g58841_da
ec0/g58841_db
ec0/g58841_sb
ec0/n_7723
ec0/n_7332
ec0/g58826_sb
ec0/n_4101
ec0/g63587_da
ec0/g63587_sb
ec0/g57096_db
ec0/g57896_sb
ec0/g57896_db
ec0/g57069_db
ec0/n_10699
ec0/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__1__Q
ec0/n_10895
ec0/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__35__Q
ec0/n_8968
ec0/n_11731
ec0/n_10705
ec0/n_10891
ec0/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__36__Q
ec0/g58019_da
ec0/g58019_sb
ec0/g57900_sb
ec0/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__0__Q
ec0/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__0__Q
ec0/g57139_db
ec0/g58008_db
ec0/n_9786
ec0/n_11702
ec0/n_8945
ec0/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_11__465
ec0/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__36__Q
ec0/n_11336
ec0/g58284_da
ec0/g58284_db
ec0/g58574_da
ec0/g58574_sb
ec0/n_9194
ec0/g58574_db
ec0/n_8952
ec0/n_9773
ec0/g58018_da
ec0/g58018_db
ec0/g57149_da
ec0/g57167_sb
ec0/g64928_da
ec0/g64928_sb
ec0/n_4315
ec0/g65065_da
ec0/g62355_da
ec0/g62355_sb
ec0/g62355_db
ec0/g62421_da
ec0/g62421_db
ec0/n_6009
ec0/g62936_da
ec0/g62936_db
ec0/g65415_sb
ec0/n_12015
ec0/n_13693
ec0/n_11938
ec0/n_3514
ec0/g65413_da
ec0/g65413_db
ec0/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__5__Q
ec0/g62515_da
ec0/g62515_sb
ec0/n_6395
ec0/g65049_db
ec0/n_4322
ec0/g65049_da
ec0/n_6485
ec0/g62541_da
ec0/g62541_db
ec0/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__2__Q
ec0/n_12508
ec0/n_12120
ec0/n_12082
ec0/g62358_sb
ec0/g62358_da
ec0/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__2__Q
ec0/n_12911
ec0/g65414_sb
ec0/n_12688
ec0/n_5950
ec0/g60672_db
ec0/g67489_p
ec0/g65522_p1
ec0/n_1175
ec0/n_1416
ec0/wishbone_slave_unit_pci_initiator_sm_latency_timer_3_
ec0/n_1011
ec0/n_1226
ec0/g65510_p
ec0/n_1178
ec0/g67514_p
ec0/n_1658
ec0/n_4663
ec0/g60671_db
ec0/g60671_da
ec0/n_5630
ec0/g62080_db
ec0/configuration_wb_err_data_580
ec0/g62098_db
ec0/n_5606
ec0/configuration_wb_err_data_571
ec0/n_7471
ec0/n_5576
ec0/g62120_db
ec0/configuration_wb_err_data_577
ec0/n_2849
ec0/n_2848
ec0/n_544
ec0/g65808_p
ec0/g65808_AP
ec0/g65808_BP
ec0/n_7212
ec0/n_1105
ec0/g61843_da
ec0/n_1978
ec0/g61831_da
ec0/n_4122
ec0/g61831_sb
ec0/g63533_da
ec0/g63533_db
ec0/g59796_da
ec0/wishbone_slave_unit_pci_initiator_if_intermediate_be_reg_1__Q
ec0/n_7621
ec0/g53893_db
ec0/n_13541
ec0/g59799_da
ec0/g54164_sb
ec0/g54166_da
ec0/g54166_sb
ec0/g54170_sb
ec0/g54170_da
ec0/wishbone_slave_unit_pcim_if_wbw_cbe_in_417
ec0/g66945_p
ec0/wishbone_slave_unit_fifos_wbr_be_in
ec0/wbu_sel_in
ec0/g58826_da
ec0/wishbone_slave_unit_wishbone_slave_d_incoming_reg_32__Q
ec0/n_8615
ec0/g58826_db
ec0/FE_OFN196_n_9230
ec0/n_9230
ec0/g57096_da
ec0/n_9139
ec0/g57096_sb
ec0/g57896_da
ec0/n_11672
ec0/FE_RN_397_0
ec0/FE_RN_398_0
ec0/n_12567
ec0/n_11727
ec0/n_9924
ec0/n_8914
ec0/g57150_sb
ec0/n_9771
ec0/g58019_db
ec0/n_9225
ec0/g57900_da
ec0/g57900_db
ec0/n_11610
ec0/g57139_da
ec0/g57977_sb
ec0/FE_OFN518_n_9823
ec0/g57139_sb
ec0/n_8485
ec0/n_8550
ec0/g58606_sb
ec0/g58271_sb
ec0/g58271_da
ec0/g57408_da
ec0/g57408_db
ec0/n_11316
ec0/g57421_db
ec0/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__21__Q
ec0/g58018_sb
ec0/g57149_db
ec0/g65065_sb
ec0/n_11839
ec0/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__20__Q
ec0/n_11800
ec0/n_6889
ec0/g62421_sb
ec0/n_3709
ec0/n_3513
ec0/g65415_da
ec0/g65415_db
ec0/g52528_sb
ec0/g52528_da
ec0/g65413_sb
ec0/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__15__Q
ec0/g63174_db
ec0/n_6548
ec0/g62515_db
ec0/g62579_da
ec0/g62579_sb
ec0/g62579_db
ec0/g64895_db
ec0/n_3698
ec0/g64895_da
ec0/g65049_sb
ec0/n_4502
ec0/g64751_da
ec0/g64751_db
ec0/g64762_sb
ec0/g64762_db
ec0/n_6883
ec0/g62358_db
ec0/n_13057
ec0/g62763_sb
ec0/g62763_da
ec0/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__36__Q
ec0/g65414_da
ec0/n_4230
ec0/g65414_db
ec0/g62966_db
ec0/n_6985
ec0/g60672_da
ec0/g60682_sb
ec0/wbu_latency_tim_val_in_246
ec0/n_560
ec0/n_561
ec0/n_1417
ec0/n_1714
ec0/wishbone_slave_unit_pci_initiator_sm_latency_timer_0_
ec0/wishbone_slave_unit_pci_initiator_sm_latency_timer_1_
ec0/n_3447
ec0/n_6982
ec0/n_4825
ec0/n_3059
ec0/n_5631
ec0/g62079_db
ec0/configuration_wb_err_addr_539
ec0/n_5555
ec0/g62138_db
ec0/g54039_sb
ec0/n_5231
ec0/g62074_db
ec0/g62073_da
ec0/g62073_sb
ec0/conf_wb_err_bc_in_846
ec0/n_832
ec0/n_715
ec0/n_8529
ec0/n_7315
ec0/n_5642
ec0/n_13750
ec0/n_13553
ec0/g61831_db
ec0/g65269_da
ec0/g65269_db
ec0/g53893_da
ec0/g53893_sb
ec0/n_13229
ec0/g54164_da
ec0/g53900_db
ec0/g54170_db
ec0/n_4104
ec0/g63584_db
ec0/n_12829
ec0/g57957_da
ec0/g57957_sb
ec0/g57957_db
ec0/g57069_da
ec0/n_9866
ec0/g57069_sb
ec0/g57946_db
ec0/g57946_da
ec0/FE_RN_197_0
ec0/n_11707
ec0/n_8890
ec0/g58588_db
ec0/n_1800
ec0/g57150_da
ec0/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__1__Q
ec0/g57150_db
ec0/g57164_sb
ec0/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__32__Q
ec0/n_11641
ec0/g57977_db
ec0/n_9824
ec0/g57977_da
ec0/g57436_sb
ec0/n_9509
ec0/g58299_da
ec0/n_10622
ec0/g58298_db
ec0/g58271_db
ec0/n_9530
ec0/g57408_sb
ec0/g58284_sb
ec0/n_11738
ec0/n_10947
ec0/n_12442
ec0/g67142_p
ec0/n_1287
ec0/n_10918
ec0/FE_RN_101_0
ec0/g57987_da
ec0/g57987_sb
ec0/n_12742
ec0/n_12336
ec0/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__15__Q
ec0/n_12604
ec0/g64923_sb
ec0/g62499_db
ec0/n_3723
ec0/g64878_db
ec0/g64849_da
ec0/g64849_sb
ec0/g64878_da
ec0/g64878_sb
ec0/g62409_sb
ec0/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__22__Q
ec0/g52528_db
ec0/wbs_wbb3_2_wbb2_dat_o_i_102
ec0/g63174_da
ec0/g63174_sb
ec0/n_12189
ec0/n_5796
ec0/g64985_db
ec0/n_3648
ec0/FE_OFN592_n_4490
ec0/g64895_sb
ec0/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__36__Q
ec0/n_6121
ec0/g64751_sb
ec0/n_13118
ec0/g62972_sb
ec0/g64762_da
ec0/n_4491
ec0/n_6117
ec0/g62763_db
ec0/n_1959
ec0/g59377_p
ec0/wishbone_slave_unit_pci_initiator_sm_latency_timer_7_
ec0/n_1716
ec0/g60672_sb
ec0/n_1715
ec0/wishbone_slave_unit_pci_initiator_sm_latency_timer_6_
ec0/g60321_p
ec0/n_2034
ec0/n_1098
ec0/n_3446
ec0/n_4664
ec0/g60674_db
ec0/n_4659
ec0/g60690_da
ec0/g60690_db
ec0/n_3041
ec0/n_2818
ec0/n_3051
ec0/n_5609
ec0/g62095_db
ec0/n_2626
ec0/n_5566
ec0/g62130_db
ec0/n_5601
ec0/g62101_db
ec0/n_2846
ec0/FE_OFN1097_n_5592
ec0/n_4811
ec0/configuration_wb_err_addr
ec0/n_5718
ec0/g62126_db
ec0/configuration_wb_err_addr_557
ec0/n_5570
ec0/n_5637
ec0/g62074_da
ec0/g62141_sb
ec0/g62074_sb
ec0/g67048_db
ec0/g67360_p
ec0/n_6942
ec0/n_1112
ec0/n_1202
ec0/n_14387
ec0/n_13753
ec0/n_13555
ec0/g53945_da
ec0/n_13499
ec0/g53945_db
ec0/g65269_sb
ec0/n_13491
ec0/n_13327
ec0/g54164_db
ec0/wishbone_slave_unit_pci_initiator_if_intermediate_be_reg_3__Q
ec0/n_13543
ec0/g53900_da
ec0/n_213
ec0/g58838_sb
ec0/g58838_da
ec0/g58838_db
ec0/n_8676
ec0/n_4102
ec0/g63586_db
ec0/g63586_da
ec0/g63584_da
ec0/g63585_sb
ec0/n_9848
ec0/g57080_sb
ec0/g57080_da
ec0/g57080_db
ec0/n_11662
ec0/g57946_sb
ec0/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__1__Q
ec0/n_11466
ec0/g58588_sb
ec0/g58588_da
ec0/n_8560
ec0/n_11600
ec0/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__1__Q
ec0/g57164_da
ec0/g57164_db
ec0/g57104_db
ec0/g57104_da
ec0/g57104_sb
ec0/n_10579
ec0/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__35__Q
ec0/g57436_db
ec0/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__35__Q
ec0/g57436_da
ec0/g58296_db
ec0/g58299_sb
ec0/g58296_sb
ec0/g58296_da
ec0/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__32__Q
ec0/g58298_sb
ec0/g58298_da
ec0/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__34__Q
ec0/n_9030
ec0/g57435_sb
ec0/g57435_da
ec0/g58293_sb
ec0/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__21__Q
ec0/FE_OFN1711_n_9320
ec0/g58251_sb
ec0/g58251_da
ec0/n_9810
ec0/g57987_db
ec0/n_6305
ec0/g62625_da
ec0/g62625_db
ec0/g64923_db
ec0/n_3682
ec0/g64923_da
ec0/n_6585
ec0/g62499_da
ec0/g64849_db
ec0/n_6781
ec0/g62409_da
ec0/g62409_db
ec0/g64794_db
ec0/n_12863
ec0/n_12605
ec0/n_12795
ec0/FE_RN_212_0
ec0/g64985_da
ec0/g64985_sb
ec0/g62758_db
ec0/n_2029
ec0/g65669_sb
ec0/g65669_da
ec0/g62760_sb
ec0/g62760_da
ec0/g62760_db
ec0/g62972_db
ec0/n_1849
ec0/n_5938
ec0/g62972_da
ec0/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__36__Q
ec0/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__36__Q
ec0/n_5800
ec0/n_12248
ec0/g65670_db
ec0/g65670_da
ec0/g65670_sb
ec0/n_2559
ec0/g59092_sb
ec0/n_104
ec0/g63989_p
ec0/n_2262
ec0/n_2218
ec0/n_247
ec0/n_3455
ec0/n_4202
ec0/n_6984
ec0/g60674_da
ec0/n_3227
ec0/g60671_sb
ec0/g60690_sb
ec0/FE_OCPN1969_n_15445
ec0/n_7220
ec0/configuration_sync_isr_2_meta_bckp_bit
ec0/configuration_sync_isr_2_sync_del_bit
ec0/configuration_sync_isr_2_delayed_del_bit_reg_Q
ec0/configuration_sync_isr_2_delayed_del_bit
ec0/n_5232
ec0/g54040_sb
ec0/g62107_sb
ec0/g62107_da
ec0/n_5593
ec0/g62107_db
ec0/n_5552
ec0/g62141_da
ec0/g62141_db
ec0/g67048_da
ec0/g67048_sb
ec0/n_13824
ec0/n_13692
ec0/n_6940
ec0/n_14392
ec0/n_13494
ec0/wishbone_slave_unit_pci_initiator_if_intermediate_be_reg_0__Q
ec0/g54158_db
ec0/n_13689
ec0/g54158_sb
ec0/g54160_sb
ec0/g53900_sb
ec0/g54160_db
ec0/n_294
ec0/g58828_db
ec0/g58828_da
ec0/wishbone_slave_unit_wishbone_slave_d_incoming_reg_34__Q
ec0/g58828_sb
ec0/n_14391
ec0/g63586_sb
ec0/g63584_sb
ec0/g58179_da
ec0/g58179_sb
ec0/g58179_db
ec0/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__1__Q
ec0/n_10777
ec0/n_10702
ec0/g57287_db
ec0/g57287_da
ec0/g58414_sb
ec0/n_10903
ec0/FE_OCPN1996_FE_OFN1711_n_9320
ec0/n_10880
ec0/n_11720
ec0/n_12564
ec0/g57988_da
ec0/g57988_sb
ec0/n_10838
ec0/n_10882
ec0/FE_RN_195_0
ec0/FE_RN_196_0
ec0/n_11726
ec0/n_11300
ec0/g57433_sb
ec0/n_9217
ec0/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__34__Q
ec0/g57435_db
ec0/n_10357
ec0/n_9031
ec0/g58293_da
ec0/g58293_db
ec0/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__2__Q
ec0/g57430_db
ec0/n_10359
ec0/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__2__Q
ec0/g58251_db
ec0/n_9043
ec0/g57113_da
ec0/g57113_sb
ec0/n_12939
ec0/n_12743
ec0/g62625_sb
ec0/g62890_sb
ec0/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__20__Q
ec0/n_12308
ec0/n_12034
ec0/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__20__Q
ec0/n_3760
ec0/g64794_da
ec0/g64794_sb
ec0/n_11889
ec0/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__15__Q
ec0/g65070_da
ec0/g65070_sb
ec0/n_12778
ec0/n_6123
ec0/g62758_da
ec0/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__36__Q
ec0/g62758_sb
ec0/g65669_db
ec0/g65672_db
ec0/n_2455
ec0/g65672_da
ec0/g65931_da
ec0/g65931_db
ec0/g63171_da
ec0/g63171_sb
ec0/g63171_db
ec0/n_2181
ec0/g63164_sb
ec0/g63164_da
ec0/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__36__Q
ec0/g65883_da
ec0/g65883_sb
ec0/g59092_da
ec0/n_3495
ec0/g59092_db
ec0/n_3443
ec0/n_4660
ec0/n_4858
ec0/n_7031
ec0/n_5748
ec0/g59226_db
ec0/n_4691
ec0/n_2906
ec0/n_4167
ec0/wbu_latency_tim_val_in_244
ec0/wbu_latency_tim_val_in
ec0/n_4899
ec0/n_3043
ec0/FE_OCPN1967_n_15445
ec0/pci_resi_conf_soft_res_in
ec0/configuration_sync_isr_2_sync_bckp_bit
ec0/configuration_sync_isr_2_meta_del_bit
ec0/n_925
ec0/configuration_set_isr_bit2
ec0/configuration_set_isr_bit2_reg_Q
ec0/n_5730
ec0/n_4883
ec0/n_3109
ec0/configuration_icr_bit_2967
ec0/n_4144
ec0/configuration_wb_err_data_576
ec0/n_5638
ec0/g62073_db
ec0/g62075_db
ec0/g62075_sb
ec0/n_8531
ec0/g59093_da
ec0/g59093_db
ec0/n_716
ec0/g59093_sb
ec0/g52877_sb
ec0/n_13826
ec0/g63315_p
ec0/wishbone_slave_unit_pci_initiator_if_posted_write_req
ec0/n_13550
ec0/n_13329
ec0/n_13548
ec0/n_13233
ec0/g54158_da
ec0/wishbone_slave_unit_pcim_if_wbw_cbe_in
ec0/g54160_da
ec0/g54168_sb
ec0/g54168_da
ec0/g52880_db
ec0/g59097_db
ec0/FE_OFN1335_n_9372
ec0/n_8611
ec0/g52880_da
ec0/g52879_da
ec0/g52879_sb
ec0/g52880_sb
ec0/n_8530
ec0/g59097_da
ec0/n_8782
ec0/n_9608
ec0/n_11433
ec0/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__0__Q
ec0/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__0__Q
ec0/g58149_db
ec0/FE_OFN500_n_9697
ec0/n_9643
ec0/g57287_sb
ec0/n_9000
ec0/g58414_da
ec0/g58414_db
ec0/g57557_da
ec0/g57557_sb
ec0/g57114_sb
ec0/g57114_da
ec0/n_9808
ec0/g57988_db
ec0/n_8947
ec0/n_11712
ec0/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__35__Q
ec0/g57433_db
ec0/g57433_da
ec0/n_10823
ec0/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__4__Q
ec0/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__4__Q
ec0/g57430_sb
ec0/g57430_da
ec0/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__30__Q
ec0/g58242_da
ec0/g58242_sb
ec0/g57394_db
ec0/g57394_da
ec0/g57394_sb
ec0/g57113_db
ec0/g65398_da
ec0/g65398_sb
ec0/n_6097
ec0/g62890_da
ec0/g62890_db
ec0/n_1576
ec0/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__36__Q
ec0/g62499_sb
ec0/FE_OFN1154_n_6391
ec0/n_6433
ec0/g65050_db
ec0/g65050_sb
ec0/n_6156
ec0/g65070_db
ec0/n_3606
ec0/g62701_db
ec0/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__15__Q
ec0/n_5924
ec0/n_13136
ec0/n_11958
ec0/g65672_sb
ec0/FE_OFN1145_n_6391
ec0/g65931_sb
ec0/FE_OFN1142_n_6391
ec0/FE_OFN364_n_6391
ec0/n_12379
ec0/n_11961
ec0/g65879_da
ec0/g65879_sb
ec0/g65879_db
ec0/n_5808
ec0/g63164_db
ec0/n_1575
ec0/g65883_db
ec0/g58611_db
ec0/n_5713
ec0/g60603_db
ec0/g60603_sb
ec0/n_4857
ec0/g59226_da
ec0/n_5728
ec0/wbu_latency_tim_val_in_245
ec0/g59226_sb
ec0/n_2819
ec0/n_2839
ec0/n_2823
ec0/FE_OCPN1966_n_15445
ec0/configuration_sync_isr_2_delayed_bckp_bit_reg_Q
ec0/n_8432
ec0/n_7571
ec0/configuration_sync_isr_2_delayed_bckp_bit
ec0/configuration_sync_isr_2_del_bit_reg_Q
ec0/n_1084
ec0/n_72
ec0/n_3247
ec0/g62076_sb
ec0/g62076_da
ec0/n_5636
ec0/g62075_da
ec0/n_14396
ec0/g52877_da
ec0/g52877_db
ec0/g52876_db
ec0/g52876_sb
ec0/g52876_da
ec0/g59239_sb
ec0/n_7028
ec0/n_4719
ec0/g53898_da
ec0/g53898_sb
ec0/g53891_da
ec0/g53891_db
ec0/g53891_sb
ec0/n_13227
ec0/n_15978
ec0/g59799_db
ec0/wishbone_slave_unit_del_sync_bc_out_reg_1__Q
ec0/g54168_db
ec0/n_526
ec0/n_211
ec0/g52879_db
ec0/wishbone_slave_unit_pcim_if_del_bc_in_382
ec0/wishbone_slave_unit_del_sync_bc_out_reg_2__Q
ec0/n_12832
ec0/n_14393
ec0/g59097_sb
ec0/FE_OFN200_n_9140
ec0/n_9140
ec0/n_16439
ec0/g57318_sb
ec0/g58169_sb
ec0/g57318_da
ec0/g57318_db
ec0/g58138_db
ec0/g58138_sb
ec0/g58149_da
ec0/g58149_sb
ec0/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__34__Q
ec0/n_10300
ec0/g57557_db
ec0/FE_RN_155_0
ec0/n_10907
ec0/FE_RN_153_0
ec0/FE_RN_154_0
ec0/n_11632
ec0/g57114_db
ec0/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__32__Q
ec0/g57129_db
ec0/n_11733
ec0/n_9918
ec0/n_8961
ec0/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__32__Q
ec0/g58301_sb
ec0/g57438_db
ec0/n_10355
ec0/FE_OFN1256_n_8567
ec0/g58242_db
ec0/n_9549
ec0/n_10374
ec0/g57152_sb
ec0/g57152_da
ec0/g57152_db
ec0/n_10109
ec0/n_6081
ec0/n_3520
ec0/g65398_db
ec0/g65873_da
ec0/g65873_db
ec0/n_12117
ec0/FE_OCPN1893_FE_OFN1474_n_14995
ec0/g62607_sb
ec0/n_6338
ec0/g62607_da
ec0/g62607_db
ec0/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__2__Q
ec0/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__236
ec0/g62563_da
ec0/g62563_sb
ec0/g62563_db
ec0/n_3620
ec0/g65050_da
ec0/g62701_da
ec0/g62701_sb
ec0/g62979_sb
ec0/g62979_da
ec0/g62979_db
ec0/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__15__Q
ec0/n_6372
ec0/g62590_da
ec0/g62590_db
ec0/n_3691
ec0/g62590_sb
ec0/n_11959
ec0/g62611_sb
ec0/n_12501
ec0/g63006_sb
ec0/g63006_da
ec0/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__3__Q
ec0/n_5870
ec0/n_12904
ec0/n_11962
ec0/g62754_sb
ec0/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__36__Q
ec0/n_6129
ec0/g63159_sb
ec0/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__3__Q
ec0/n_5819
ec0/n_4892
ec0/n_7602
ec0/g60603_da
ec0/wbu_latency_tim_val_in_248
ec0/n_15731
ec0/n_16429
ec0/n_15606
ec0/wbu_latency_tim_val_in_243
ec0/g60674_sb
ec0/n_7607
ec0/n_2845
ec0/n_4852
ec0/n_4648
ec0/n_3056
ec0/configuration_isr_bit_1457
ec0/configuration_isr_bit_618
ec0/n_4146
ec0/n_3117
ec0/n_3245
ec0/configuration_icr_bit_2961
ec0/n_7817
ec0/n_7819
ec0/n_4780
ec0/g62076_db
ec0/n_5635
ec0/g62077_sb
ec0/FE_RN_165_0
ec0/n_14397
ec0/g52878_sb
ec0/g52878_da
ec0/g59239_da
ec0/n_7714
ec0/g59239_db
ec0/n_7077
ec0/g53898_db
ec0/g63338_p
ec0/n_15054
ec0/n_2354
ec0/wishbone_slave_unit_pci_initiator_if_write_req_int
ec0/g59763_sb
ec0/g59763_da
ec0/g52881_db
ec0/wishbone_slave_unit_pcim_if_del_bc_in_383
ec0/n_8598
ec0/wishbone_slave_unit_pcim_if_del_bc_in
ec0/n_8723
ec0/n_8597
ec0/g57308_sb
ec0/g57308_da
ec0/n_9622
ec0/g58169_da
ec0/g58169_db
ec0/g57276_sb
ec0/g57276_da
ec0/n_9658
ec0/g58138_da
ec0/g57276_db
ec0/n_10898
ec0/n_9922
ec0/n_8967
ec0/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__35__Q
ec0/g57555_sb
ec0/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__34__Q
ec0/n_10908
ec0/FE_RN_93_0
ec0/g57552_db
ec0/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__32__Q
ec0/g57552_sb
ec0/n_10841
ec0/g57129_da
ec0/n_9227
ec0/g57129_sb
ec0/n_8965
ec0/n_8943
ec0/n_9910
ec0/n_1822
ec0/n_8957
ec0/g58301_db
ec0/g58301_da
ec0/g57438_da
ec0/n_9029
ec0/g57438_sb
ec0/g58294_db
ec0/g58294_sb
ec0/g57385_db
ec0/g57385_sb
ec0/g57385_da
ec0/n_9768
ec0/g58021_da
ec0/g58021_db
ec0/g62898_da
ec0/g62898_db
ec0/g62898_sb
ec0/g65889_sb
ec0/g65873_sb
ec0/n_4400
ec0/n_4399
ec0/g64912_db
ec0/n_12457
ec0/g65028_da
ec0/g65028_sb
ec0/g62994_sb
ec0/g62994_da
ec0/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__2__Q
ec0/n_4156
ec0/n_12446
ec0/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__249
ec0/n_3692
ec0/g62611_da
ec0/n_3738
ec0/FE_OFN320_g66077_p
ec0/n_12677
ec0/g63006_db
ec0/n_3571
ec0/g65309_sb
ec0/n_13034
ec0/n_12814
ec0/n_12246
ec0/n_11819
ec0/n_11960
ec0/g62761_da
ec0/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__36__Q
ec0/g62761_sb
ec0/g62754_da
ec0/g62754_db
ec0/g63159_da
ec0/g63159_db
ec0/g58611_da
ec0/g58611_sb
ec0/n_7601
ec0/n_7459
ec0/n_7461
ec0/n_15732
ec0/n_15733
ec0/g63362_p
ec0/n_7604
ec0/n_2797
ec0/n_7606
ec0/n_7605
ec0/n_7465
ec0/n_7469
ec0/n_2912
ec0/n_15627
ec0/n_4855
ec0/configuration_pci_err_addr_479
ec0/n_3180
ec0/configuration_isr_bit_1461
ec0/n_536
ec0/n_3799
ec0/configuration_isr_bit_2975
ec0/n_8508
ec0/n_7742
ec0/n_369
ec0/n_7472
ec0/n_7473
ec0/n_7474
ec0/n_5634
ec0/g62077_da
ec0/g62077_db
ec0/FE_RN_166_0
ec0/FE_RN_167_0
ec0/g52878_db
ec0/n_14394
ec0/g63206_p
ec0/n_416
ec0/n_1659
ec0/n_5228
ec0/g61617_p
ec0/wishbone_slave_unit_pci_initiator_if_read_count_3_
ec0/wishbone_slave_unit_pci_initiator_if_read_count_reg_3__Q
ec0/n_7544
ec0/g17_p
ec0/n_2355
ec0/n_1780
ec0/g59763_db
ec0/n_2328
ec0/n_7625
ec0/wishbone_slave_unit_del_sync_bc_out_reg_0__Q
ec0/wishbone_slave_unit_del_sync_bc_out_reg_3__Q
ec0/n_8796
ec0/n_14388
ec0/g52881_da
ec0/g52881_sb
ec0/n_11442
ec0/g57308_db
ec0/n_8966
ec0/n_11478
ec0/n_11706
ec0/n_8889
ec0/g58412_da
ec0/g58412_sb
ec0/n_9205
ec0/g58412_db
ec0/g57555_da
ec0/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__32__Q
ec0/n_10810
ec0/g57552_da
ec0/n_9207
ec0/g58410_da
ec0/g58410_db
ec0/g58410_sb
ec0/g57897_db
ec0/g57897_da
ec0/n_11700
ec0/n_8553
ec0/g58595_db
ec0/g57598_db
ec0/n_10285
ec0/n_9511
ec0/g58294_da
ec0/g57431_da
ec0/g57431_sb
ec0/g57431_db
ec0/n_11359
ec0/g58256_sb
ec0/g58021_sb
ec0/g57990_sb
ec0/g57990_da
ec0/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__21__Q
ec0/n_1860
ec0/g65889_da
ec0/g65889_db
ec0/FE_OCPN1892_FE_OFN1474_n_14995
ec0/n_12122
ec0/g63153_db
ec0/n_1861
ec0/g65888_sb
ec0/g64912_da
ec0/g64912_sb
ec0/g65432_db
ec0/n_4337
ec0/g65028_db
ec0/g62416_db
ec0/n_5894
ec0/g62994_db
ec0/g65395_da
ec0/g65395_db
ec0/g65395_sb
ec0/g64892_sb
ec0/g64892_da
ec0/g64903_db
ec0/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__237
ec0/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__3__Q
ec0/n_6334
ec0/g62611_db
ec0/g64819_db
ec0/n_3740
ec0/g64819_da
ec0/g65309_da
ec0/n_12236
ec0/g65673_db
ec0/n_6119
ec0/g62761_db
ec0/g65668_db
ec0/n_3548
ec0/g65340_da
ec0/g65340_sb
ec0/g65340_db
ec0/wbu_latency_tim_val_in_249
ec0/n_7467
ec0/n_7600
ec0/n_2905
ec0/n_4641
ec0/n_3037
ec0/n_7463
ec0/n_7468
ec0/n_2969
ec0/n_4125
ec0/n_5701
ec0/configuration_wb_err_cs_bit9
ec0/n_6218
ec0/n_535
ec0/n_1120
ec0/n_3800
ec0/configuration_command_bit
ec0/n_3235
ec0/n_4088
ec0/n_2847
ec0/configuration_pci_err_data_507
ec0/g62072_sb
ec0/g59390_p
ec0/n_4703
ec0/FE_RN_169_0
ec0/g59129_p
ec0/wishbone_slave_unit_pci_initiator_if_read_count_2_
ec0/n_7333
ec0/n_660
ec0/n_2014
ec0/n_7079
ec0/n_15262
ec0/g65573_p
ec0/n_2801
ec0/n_2088
ec0/g67709_p
ec0/n_8677
ec0/n_8680
ec0/n_8596
ec0/wishbone_slave_unit_wishbone_slave_map
ec0/n_1323
ec0/wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg_Q
ec0/n_9920
ec0/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__35__Q
ec0/g58104_sb
ec0/n_10806
ec0/g57555_db
ec0/g58262_sb
ec0/g57899_db
ec0/g57899_sb
ec0/g57897_sb
ec0/g58446_da
ec0/g58446_sb
ec0/g58595_sb
ec0/g58595_da
ec0/g57596_db
ec0/n_9038
ec0/g58263_da
ec0/g58263_db
ec0/g57598_da
ec0/n_11303
ec0/g58256_da
ec0/n_9040
ec0/g58256_db
ec0/g58576_sb
ec0/g57990_db
ec0/FE_RN_100_0
ec0/n_10041
ec0/n_12375
ec0/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__36__Q
ec0/n_5836
ec0/g63153_da
ec0/g65888_db
ec0/g65888_da
ec0/n_5997
ec0/g62942_da
ec0/g62942_db
ec0/n_4673
ec0/g65432_da
ec0/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__2__Q
ec0/g65432_sb
ec0/g62416_da
ec0/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__2__Q
ec0/g62416_sb
ec0/n_6766
ec0/n_4245
ec0/g65383_da
ec0/g65383_sb
ec0/g62573_db
ec0/n_4412
ec0/g64892_db
ec0/g64903_sb
ec0/g64903_da
ec0/n_12454
ec0/g64819_sb
ec0/g65309_db
ec0/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__36__Q
ec0/n_13319
ec0/n_12960
ec0/n_1958
ec0/g65673_da
ec0/n_12667
ec0/n_11949
ec0/g65098_sb
ec0/n_1960
ec0/g65668_da
ec0/g64955_sb
ec0/n_7599
ec0/n_14917
ec0/n_7261
ec0/n_7457
ec0/g66446_p
ec0/n_231
ec0/n_14911
ec0/n_7237
ec0/n_4683
ec0/configuration_pci_err_addr_480
ec0/n_4849
ec0/n_4813
ec0/configuration_icr_bit2_0
ec0/configuration_isr_bit_631
ec0/n_2898
ec0/n_7820
ec0/g64632_p
ec0/n_15435
ec0/configuration_pci_err_addr
ec0/n_8477
ec0/n_7610
ec0/n_8474
ec0/n_7612
ec0/g67156_p
ec0/FE_RN_168_0
ec0/FE_RN_170_0
ec0/n_1660
ec0/n_4859
ec0/n_5229
ec0/g60409_sb
ec0/g63925_p
ec0/FE_RN_237_0
ec0/g63530_db
ec0/g63530_sb
ec0/g63530_da
ec0/wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_36__Q
ec0/g58837_da
ec0/g58837_sb
ec0/g58837_db
ec0/n_1721
ec0/wishbone_slave_unit_wishbone_slave_mrl_en_reg_Q
ec0/n_7542
ec0/n_12828
ec0/n_11705
ec0/n_8888
ec0/g58164_da
ec0/g58164_sb
ec0/g58164_db
ec0/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__4__Q
ec0/g58104_da
ec0/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__4__Q
ec0/n_10576
ec0/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__36__Q
ec0/FE_RN_94_0
ec0/FE_RN_95_0
ec0/n_9039
ec0/g58262_da
ec0/g58262_db
ec0/n_10890
ec0/n_9138
ec0/g57899_da
ec0/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__30__Q
ec0/n_10561
ec0/n_9199
ec0/g58446_db
ec0/n_10797
ec0/g57596_da
ec0/g58263_sb
ec0/g57598_sb
ec0/n_10372
ec0/n_11451
ec0/g58161_db
ec0/g57400_sb
ec0/g57400_da
ec0/g57400_db
ec0/g57118_sb
ec0/n_9805
ec0/g57118_da
ec0/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__2__Q
ec0/g64870_da
ec0/g64870_sb
ec0/n_12676
ec0/n_12376
ec0/g63153_sb
ec0/g62991_da
ec0/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__27__Q
ec0/g62991_sb
ec0/g62942_sb
ec0/n_12263
ec0/n_11978
ec0/g65383_db
ec0/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__2__Q
ec0/n_6407
ec0/g62573_da
ec0/g62998_sb
ec0/n_12790
ec0/g64991_sb
ec0/g64991_da
ec0/g65897_sb
ec0/g65897_da
ec0/g62997_sb
ec0/g62997_da
ec0/g65673_sb
ec0/n_13053
ec0/g65098_da
ec0/g62363_db
ec0/n_3595
ec0/g65668_sb
ec0/g64955_da
ec0/n_3663
ec0/g64955_db
ec0/n_14915
ec0/n_7263
ec0/n_7455
ec0/n_7011
ec0/n_7009
ec0/n_15699
ec0/n_15434
ec0/n_2862
ec0/n_7452
ec0/n_7280
ec0/pciu_am1_in_520
ec0/g67536_p
ec0/n_6995
ec0/n_2824
ec0/n_2614
ec0/g60635_db
ec0/configuration_sync_pci_err_cs_8_delayed_del_bit_reg_Q
ec0/configuration_sync_pci_err_cs_8_sync_del_bit
ec0/configuration_wb_err_cs_bit8
ec0/n_8510
ec0/n_7743
ec0/n_24
ec0/n_15436
ec0/n_7475
ec0/g61572_p
ec0/n_8453
ec0/n_8454
ec0/n_7611
ec0/g61581_p
ec0/n_676
ec0/g58656_p
ec0/n_7094
ec0/n_4851
ec0/n_5646
ec0/n_703
ec0/wishbone_slave_unit_pci_initiator_if_read_count_1_
ec0/n_9
ec0/g60409_da
ec0/g60409_db
ec0/n_4591
ec0/n_3437
ec0/n_21
ec0/n_3429
ec0/FE_RN_238_0
ec0/FE_RN_236_0
ec0/FE_RN_235_0
ec0/FE_RN_244_0
ec0/wishbone_slave_unit_wishbone_slave_pref_en_reg_Q
ec0/n_7718
ec0/n_7719
ec0/n_5735
ec0/configuration_meta_command_bit
ec0/g57302_sb
ec0/g57302_da
ec0/n_9065
ec0/g57302_db
ec0/g57334_sb
ec0/g57334_da
ec0/n_9079
ec0/g58104_db
ec0/g57334_db
ec0/n_8912
ec0/n_1821
ec0/g57554_db
ec0/g57554_da
ec0/g57554_sb
ec0/g57131_db
ec0/g57131_da
ec0/g57131_sb
ec0/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__36__Q
ec0/g57596_sb
ec0/n_1820
ec0/g58254_sb
ec0/g58254_da
ec0/n_9042
ec0/g58254_db
ec0/g57398_da
ec0/g57398_db
ec0/g57300_da
ec0/g57300_db
ec0/n_9627
ec0/g57300_sb
ec0/g58161_da
ec0/g58161_sb
ec0/n_10368
ec0/g57118_db
ec0/n_11628
ec0/g57998_db
ec0/n_4424
ec0/g64870_db
ec0/n_11992
ec0/n_12393
ec0/n_5900
ec0/g62991_db
ec0/g65357_db
ec0/n_4256
ec0/g64966_sb
ec0/n_12692
ec0/FE_RN_210_0
ec0/n_12913
ec0/g65015_sb
ec0/g65015_da
ec0/g62493_db
ec0/n_3635
ec0/FE_RN_211_0
ec0/g62573_sb
ec0/n_11976
ec0/n_12261
ec0/g62998_da
ec0/n_5886
ec0/g62998_db
ec0/g64991_db
ec0/g65897_db
ec0/n_5888
ec0/g62997_db
ec0/g65098_db
ec0/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__3__Q
ec0/n_6875
ec0/g62363_da
ec0/g62677_db
ec0/n_16852
ec0/n_15698
ec0/n_3308
ec0/n_14913
ec0/n_7271
ec0/g60605_db
ec0/n_15623
ec0/configuration_sync_pci_err_cs_8_delayed_del_bit
ec0/n_1191
ec0/g60345_p
ec0/n_4695
ec0/n_8445
ec0/n_7793
ec0/n_7794
ec0/n_7613
ec0/n_7590
ec0/n_7419
ec0/g60604_db
ec0/g60673_db
ec0/g60408_sb
ec0/n_4861
ec0/g60407_da
ec0/g60407_db
ec0/g60407_sb
ec0/n_4870
ec0/wishbone_slave_unit_pci_initiator_if_read_bound
ec0/n_4809
ec0/n_5737
ec0/n_5739
ec0/n_665
ec0/FE_OFN932_n_2700
ec0/n_16068
ec0/n_8525
ec0/n_16437
ec0/n_10407
ec0/n_10396
ec0/g58589_db
ec0/g58589_da
ec0/n_8559
ec0/g58589_sb
ec0/n_1540
ec0/n_10302
ec0/n_10473
ec0/g58190_db
ec0/n_8557
ec0/n_1542
ec0/g58593_db
ec0/n_8904
ec0/g58593_da
ec0/n_8555
ec0/g57398_sb
ec0/g58105_sb
ec0/g58105_da
ec0/g58105_db
ec0/g58029_sb
ec0/g58029_db
ec0/g57998_sb
ec0/g57998_da
ec0/n_6493
ec0/g62538_db
ec0/g65357_da
ec0/g62419_db
ec0/n_6759
ec0/n_6598
ec0/g62493_da
ec0/n_12912
ec0/n_12691
ec0/n_6356
ec0/n_4358
ec0/n_1718
ec0/g64874_sb
ec0/g62363_sb
ec0/g62677_da
ec0/n_14918
ec0/n_7228
ec0/n_6992
ec0/n_16853
ec0/n_15553
ec0/n_15552
ec0/n_15694
ec0/n_15695
ec0/n_15696
ec0/g67313_p
ec0/n_7014
ec0/n_7290
ec0/n_7460
ec0/n_15624
ec0/n_7434
ec0/n_7595
ec0/n_4860
ec0/g60408_da
ec0/n_2234
ec0/n_5758
ec0/n_15741
ec0/n_7300
ec0/FE_OFN936_n_2696
ec0/n_5741
ec0/FE_RN_57_0
ec0/FE_RN_259_0
ec0/g75084_p
ec0/n_7816
ec0/g75067_p
ec0/g58190_sb
ec0/g58190_da
ec0/g58591_sb
ec0/g58002_sb
ec0/g58593_sb
ec0/g57999_sb
ec0/g58029_da
ec0/g58189_sb
ec0/g58160_sb
ec0a/n_783
ec0a/n_326
ec0a/wbu_we_in
ec0a/n_2557
ec0a/g66223_p
ec0a/g59126_da
ec0a/g59126_sb
ec0a/g59126_db
ec0a/n_15417
ec0a/n_16952
ec0a/g75332_p
ec0a/n_15414
ec0a/FE_RN_317_0
ec0a/FE_RN_319_0
ec0a/n_8583
ec0a/n_16910
ec0a/g74660_p
ec0a/FE_RN_450_0
ec0a/n_16854
ec0a/wishbone_slave_unit_del_sync_comp_cycle_count_reg_9__Q
ec0a/n_8655
ec0a/wishbone_slave_unit_del_sync_comp_cycle_count_9_
ec0a/wbs_rty_o_1308
ec0a/n_15418
ec0a/n_15416
ec0a/FE_OCPUNCON2097_n_8660
ec0a/FE_OCPUNCON2096_n_8660
ec0a/wishbone_slave_unit_del_sync_comp_cycle_count_reg_13__Q
ec0a/n_8650
ec0a/n_2422
ec0a/n_8661
ec0a/wishbone_slave_unit_del_sync_comp_cycle_count_reg_8__Q
ec0a/wishbone_slave_unit_del_sync_comp_cycle_count_reg_14__Q
ec0a/n_8649
ec0a/n_2731
ec0a/g64371_p
ec0a/n_1992
ec0a/n_1631
ec0a/wishbone_slave_unit_del_sync_comp_cycle_count_8_
ec0a/n_4800
ec0a/n_3184
ec0a/g63428_p
ec0a/n_1994
ec0a/n_2176
ec0a/g57033_p
ec0a/n_3462
ec0a/g59367_p
ec0a/n_2474
ec0a/n_1993
ec0a/n_245
ec0a/n_3073
ec0a/n_193
ec0a/wishbone_slave_unit_del_sync_req_rty_exp_clr_reg_Q
ec0a/n_3074
ec0a/wishbone_slave_unit_del_sync_comp_cycle_count_reg_15__Q
ec0a/n_2490
ec0a/n_784
ec0a/n_206
ec0a/n_785
ec0a/n_2425
ec0a/g63208_p
ec0a/n_1327
ec0a/n_3209
ec0a/g59206_p
ec0a/n_3329
ec0a/g57878_p
ec0a/wishbone_slave_unit_del_sync_comp_cycle_count_11_
ec0a/wishbone_slave_unit_del_sync_comp_cycle_count_12_
ec0a/g59785_p
ec0a/n_2965
ec0a/n_2386
ec0a/n_8648
ec0a/n_8662
ec0a/wishbone_slave_unit_del_sync_comp_cycle_count_reg_12__Q
ec0a/wishbone_slave_unit_del_sync_comp_cycle_count_reg_11__Q
ec0a/n_2996
ec0a/n_8656
ec0a/wishbone_slave_unit_del_sync_comp_cycle_count_reg_10__Q
ec0a/wishbone_slave_unit_del_sync_sync_comp_rty_exp_clr
ec0a/n_8651
ec0a/n_6975
ec0a/g61836_da
ec0a/g61836_db
ec0a/wishbone_slave_unit_del_sync_comp_rty_exp_clr_reg_Q
ec0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__1__Q
ec0a/n_5716
ec0a/g61698_da
ec0a/g61698_db
ec0a/n_4617
ec0a/g61698_sb
ec0a/n_4613
ec0a/g61836_sb
ec0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__1__Q
ec0a/g63361_p
ec0a/wishbone_slave_unit_del_sync_comp_rty_exp_clr
ec0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__1__Q
ec0a/n_6973
ec0a/g63538_db
ec0a/g63538_da
ec0a/g63538_sb
ec0a/g63543_da
ec0a/g63543_sb
ec0a/g63543_db
ec0a/g61837_da
ec0a/g61837_db
ec0a/n_14225
ec0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__1__Q
ec0a/n_6967
ec0a/g63549_da
ec0a/g63549_sb
ec0a/n_4618
ec0a/g61837_sb
ec0a/n_14223
ec0a/n_14462
ec0a/g61842_da
ec0a/g61842_db
ec0a/n_4608
ec0a/g61842_sb
ec0a/g63549_db
ec0a/n_13893
ec0a/g63537_da
ec0a/g63537_db
ec0a/n_14277
ec0a/g63043_sb
ec0a/n_14052
ec0a/g63537_sb
ec0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__35__Q
ec0a/n_5166
ec0a/g63043_da
ec0a/g63043_db
ec0a/n_3916
ec0a/g64257_da
ec0a/g64257_db
ec0a/n_6977
ec0a/g61835_da
ec0a/g61835_db
ec0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__0__Q
ec0a/n_4599
ec0a/g63563_da
ec0a/g63563_db
ec0a/g61955_sb
ec0a/n_13950
ec0a/g64257_sb
ec0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__1__Q
ec0a/n_6958
ec0a/g61835_sb
ec0a/n_4611
ec0a/g63563_sb
ec0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__0__Q
ec0a/g61955_da
ec0a/g53267_p
ec0a/g63548_sb
ec0a/g63548_da
ec0a/g61957_db
ec0a/g63545_da
ec0a/g63545_db
ec0a/n_13906
ec0a/n_6963
ec0a/g61955_db
ec0a/g63548_db
ec0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__0__Q
ec0a/n_4609
ec0a/g61841_da
ec0a/g61841_sb
ec0a/g61957_da
ec0a/n_4597
ec0a/g61957_sb
ec0a/g63545_sb
ec0a/g64340_db
ec0a/n_14302
ec0a/g61841_db
ec0a/n_6969
ec0a/g63565_da
ec0a/g63565_db
ec0a/g63170_sb
ec0a/g63170_da
ec0a/n_3838
ec0a/n_14427
ec0a/n_14248
ec0a/n_13979
ec0a/g63565_sb
ec0a/g64340_da
ec0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__35__Q
ec0a/g64340_sb
ec0a/n_14301
ec0a/g53199_p
ec0a/g53155_p
ec0a/n_14249
ec0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__1__Q
ec0a/n_6948
ec0a/n_13978
ec0a/g63170_db
ec0a/n_4953
ec0a/n_14569
ec0a/n_14480
ec0a/g61963_db
ec0a/g63566_da
ec0a/g63566_sb
ec0a/n_14481
ec0a/n_14162
ec0a/g63544_da
ec0a/g63544_db
ec0a/g63544_sb
ec0a/g61963_da
ec0a/n_4596
ec0a/g61963_sb
ec0a/g63566_db
ec0a/n_13949
ec0a/g64123_sb
ec0a/n_14426
ec0a/n_14543
ec0a/n_14510
ec0a/g53268_p
ec0a/n_5014
ec0a/n_13947
ec0a/n_5016
ec0a/g64123_da
ec0a/g64123_db
ec0a/g63139_da
ec0a/n_3815
ec0a/g63139_sb
ec0a/n_4970
ec0a/g63139_db
ec0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__6__Q
ec0a/g63121_db
ec0a/g63121_da
ec0a/g63120_da
ec0a/g63120_db
ec0a/g64365_da
ec0a/g64365_sb
ec0a/g63121_sb
ec0a/n_3850
ec0a/g63120_sb
ec0a/g64326_da
ec0b/g57267_da
ec0b/g57267_sb
ec0b/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__30__Q
ec0b/n_9873
ec0b/g57937_db
ec0b/g57057_da
ec0b/g57057_db
ec0b/n_11485
ec0b/g57267_db
ec0b/g57057_sb
ec0b/g58220_db
ec0b/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__30__Q
ec0b/n_9262
ec0b/g58220_sb
ec0b/n_9567
ec0b/g58220_da
ec0b/n_9261
ec0b/g58265_sb
ec0b/g57590_db
ec0b/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__4__Q
ec0b/g57363_sb
ec0b/g57363_da
ec0b/g58335_sb
ec0b/g57590_sb
ec0b/n_10289
ec0b/g57590_da
ec0b/g57363_db
ec0b/g58335_db
ec0b/n_9021
ec0b/g58335_da
ec0b/g57474_db
ec0b/g58062_db
ec0b/g58062_da
ec0b/n_8990
ec0b/g58454_da
ec0b/g58454_sb
ec0b/n_16851
ec0b/g58132_sb
ec0b/n_11384
ec0b/g57474_sb
ec0b/g57474_da
ec0b/g58062_sb
ec0b/g57407_sb
ec0b/g58454_db
ec0b/g57270_sb
ec0b/g58132_da
ec0b/g57940_sb
ec0b/g57940_da
ec0b/n_10308
ec0b/n_9036
ec0b/g58270_da
ec0b/g58270_sb
ec0b/n_10417
ec0b/g57270_da
ec0b/g57270_db
ec0b/n_9073
ec0b/g58132_db
ec0b/g57063_sb
ec0b/g57063_da
ec0b/n_9130
ec0b/g57940_db
ec0b/g57546_da
ec0b/g57546_db
ec0b/g58267_sb
ec0b/g58270_db
ec0b/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__4__Q
ec0b/g57063_db
ec0b/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__4__Q
ec0b/g57546_sb
ec0b/g58267_da
ec0b/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__34__Q
ec0b/n_10290
ec0b/n_10503
ec0b/n_16850
ec0b/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__34__Q
ec0b/n_9037
ec0b/g58267_db
ec0b/g57587_db
ec0b/g57587_da
ec0b/n_9982
ec0b/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__4__Q
ec0b/n_10564
ec0b/g58607_sb
ec0b/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__4__Q
ec0b/g57587_sb
ec0b/g57201_db
ec0b/n_8900
ec0b/g58607_da
ec0b/g58607_db
ec0b/n_8549
ec0b/n_8484
ec0b/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_13__543
ec0b/g58609_sb
ec0b/g58609_da
ec0b/g57905_db
ec0b/n_10445
ec0b/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__36__Q
ec0b/n_16844
ec0b/n_354
ec0b/n_393
ec0b/g58609_db
ec0b/n_9136
ec0b/g57905_da
ec0b/g57201_da
ec0b/g57201_sb
ec0b/g58594_db
ec0b/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__36__Q
ec0b/n_8902
ec0b/g57558_da
ec0b/g57905_sb
ec0b/n_8959
ec0b/g58586_da
ec0b/g58586_db
ec0b/g58586_sb
ec0b/n_8562
ec0b/g58594_sb
ec0b/g58594_da
ec0b/n_8554
ec0b/g57558_sb
ec0b/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__36__Q
ec0b/n_1806
ec0b/n_1230
ec0b/n_9993
ec0b/n_337
ec0b/g58587_da
ec0b/n_8563
ec0b/g58587_sb
ec0b/n_1493
ec0b/n_16845
ec0b/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__36__Q
ec0b/n_10577
ec0b/g57238_db
ec0b/n_8916
ec0b/g58587_db
ec0b/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__36__Q
ec0b/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__36__Q
ec0b/n_10430
ec0b/g58094_db
ec0b/g57238_da
ec0b/n_10384
ec0b/g57366_db
ec0b/g57366_da
ec0b/n_9191
ec0b/n_9082
ec0b/g57238_sb
ec0b/n_8906
ec0b/g58592_db
ec0b/g58223_db
ec0b/n_9050
ec0b/g57366_sb
ec0b/g58596_db
ec0b/g58596_da
ec0b/g58094_da
ec0b/g58094_sb
ec0b/g58592_da
ec0b/n_1814
ec0b/g58223_da
ec0b/n_1810
ec0b/n_8552
ec0b/g58596_sb
ec0b/g57503_sb
ec0b/n_8556
ec0b/g58592_sb
ec0b/g58365_sb
ec0b/g58223_sb
ec0b/g58365_db
ec0b/g57503_da
ec0b/g57503_db
ec0b/FE_OFN245_n_9116
ec0b/g57505_db
ec0b/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__32__Q
ec0b/n_10817
ec0b/g57505_da
ec0b/g58365_da
ec0b/n_9210
ec0b/FE_OFN1278_n_8567
ec0b/n_11235
ec0b/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__32__Q
ec0b/n_10845
ec0b/g57146_sb
ec0b/g57505_sb
ec0b/g58101_sb
ec0b/g58015_sb
ec0b/n_8482
ec0b/g57094_db
ec0b/g57094_da
ec0b/g57094_sb
ec0b/g57146_da
ec0b/n_9777
ec0b/n_11604
ec0b/g57146_db
ec0b/g58101_da
ec0b/g58015_da
ec0b/g58015_db
ec0b/g57894_db
ec0b/n_9231
ec0b/g57894_da
ec0b/n_9698
ec0b/g58101_db
ec0b/g57379_sb
ec0b/g57894_sb
ec0b/g57306_db
ec0b/g57306_da
ec0b/n_9556
ec0d/g52484_db
ec0d/wishbone_slave_unit_delayed_write_data_comp_wdata_out_95
ec0d/g54219_sb
ec0d/g54182_db
ec0d/g54195_db
ec0d/g54188_sb
ec0d/g63252_p
ec0d/g54233_db
ec0d/g54219_db
ec0d/wishbone_slave_unit_delayed_write_data_comp_wdata_out_94
ec0d/g58458_sb
ec0d/g54188_da
ec0d/g54142_sb
ec0d/g54233_da
ec0d/n_13172
ec0d/g54219_da
ec0d/g54182_da
ec0d/g54182_sb
ec0d/g58458_da
ec0d/n_8989
ec0d/g58458_db
ec0d/n_13202
ec0d/n_13525
ec0d/g53917_da
ec0d/g53917_db
ec0d/n_13209
ec0d/g54189_db
ec0d/g53917_sb
ec0d/n_13108
ec0d/g54232_da
ec0d/g54189_da
ec0d/g54189_sb
ec0d/g54195_sb
ec0d/g54175_db
ec0d/n_13109
ec0d/g54184_db
ec0d/g54195_da
ec0d/n_13161
ec0d/g54232_db
ec0d/g54184_da
ec0d/FE_OFN1002_n_13221
ec0d/FE_OFN1003_n_13221
ec0d/g54143_sb
ec0d/g53932_sb
ec0d/g53932_da
ec0d/wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_9__Q
ec0d/n_13513
ec0d/g53932_db
ec0d/wishbone_slave_unit_delayed_write_data_comp_wdata_out_79
ec0d/n_833
ec0d/g67032_p
ec0d/g62065_sb
ec0d/g54199_db
ec0d/n_1004
ec0d/g53935_db
ec0d/n_13218
ec0d/g53904_sb
ec0d/g54175_da
ec0d/g54175_sb
ec0d/g54184_sb
ec0d/wishbone_slave_unit_delayed_write_data_comp_wdata_out_82
ec0d/g53935_da
ec0d/n_13537
ec0d/g53904_da
ec0d/g53904_db
ec0d/wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_12__Q
ec0d/n_13183
ec0d/g54207_da
ec0d/g54207_db
ec0d/g67003_p
ec0d/g62036_sb
ec0d/g54199_da
ec0d/g54197_db
ec0d/g67021_p
ec0d/g54237_da
ec0d/g54237_db
ec0d/FE_OFN1086_n_13249
ec0d/g54136_da
ec0d/g54136_sb
ec0d/g54237_sb
ec0d/g54213_da
ec0d/g54207_sb
ec0d/g54198_db
ec0d/g54136_db
ec0d/n_13530
ec0d/g54197_da
ec0d/g53911_db
ec0d/n_13177
ec0d/g54213_db
ec0d/wishbone_slave_unit_delayed_write_data_comp_wdata_out_89
ec0d/n_13193
ec0d/g53911_da
ec0d/g53911_sb
ec0d/g54199_sb
ec0d/g54198_da
ec0d/n_13196
ec0d/g62055_sb
ec0d/g53923_sb
ec0d/g54197_sb
ec0d/g54196_da
ec0d/g54196_db
ec0d/g54224_db
ec0d/wishbone_slave_unit_delayed_write_data_comp_wdata_out_72
ec0d/g54148_db
ec0d/wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_2__Q
ec0d/g53923_da
ec0d/n_13521
ec0d/g53923_db
ec0d/n_13168
ec0d/g54224_da
ec0d/g54174_sb
ec0d/g54148_da
ec0d/g54148_sb
ec0d/g54196_sb
ec0d/n_13219
ec0d/g54174_da
ec0d/g53939_db
ec0d/wishbone_slave_unit_delayed_write_data_comp_wdata_out_77
ec0d/g54230_db
ec0d/g54198_sb
ec0d/g54185_sb
ec0d/n_13206
ec0d/g54185_da
ec0d/g62051_db
ec0d/g53930_db
ec0d/n_13163
ec0d/g54230_da
ec0d/g54227_da
ec0d/g62051_da
ec0d/wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_26__Q
ec0d/g62051_sb
ec0d/g53919_da
ec0d/g53919_sb
ec0d/n_13166
ec0d/g54227_db
ec0d/wishbone_slave_unit_delayed_write_data_comp_wdata_out_74
ec0d/g53930_sb
ec0d/n_13248
ec0d/n_13515
ec0d/g53930_da
ec0d/n_13627
ec0d/g53919_db
ec0d/g54151_da
ec0d/g54151_db
ec0d/g54151_sb
ec0d/g54144_da
ec0d/g54144_db
ec0d/g62059_sb
ec0d/g54144_sb
ec0d/g54155_sb
ec0d/g54139_sb
ec0d/g53927_db
ec0d/n_13325
ec0d/g54220_da
ec0d/g54220_db
ec0d/g54216_sb
ec0d/g54155_da
ec0d/g54155_db
ec0d/g54139_da
ec0d/g54139_db
ec0d/g54172_sb
ec0d/g54172_db
ec0d/g62046_sb
ec0d/g54172_da
ec0d/g54173_sb
ec0d/g54173_da
ec0d/g54173_db
ec0d/g54216_da
ec0f/g65022_da
ec0f/n_3631
ec0f/FE_OFN1459_n_12306
ec0f/g62690_db
ec0f/n_4915
ec0f/FE_OFN1224_n_6624
ec0f/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__37__Q
ec0f/n_7364
ec0f/n_4511
ec0f/n_4096
ec0f/g62689_db
ec0f/n_4510
ec0f/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_14__583
ec0f/n_395
ec0f/g62690_da
ec0f/n_4907
ec0f/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_7__310
ec0f/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__37__Q
ec0f/n_7374
ec0f/g62689_da
ec0f/g62689_sb
ec0f/n_7366
ec0f/n_12245
ec0f/g62690_sb
ec0f/g62618_db
ec0f/g62618_da
ec0f/FE_OFN1434_n_12042
ec0f/g62460_sb
ec0f/n_11953
ec0f/FE_OFN1230_n_6624
ec0f/n_12675
ec0f/FE_OFN1473_n_14995
ec0f/g62618_sb
ec0f/n_4908
ec0f/n_6676
ec0f/g62460_da
ec0f/g62448_da
ec0f/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__3__Q
ec0f/g62448_sb
ec0f/n_12500
ec0f/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__5__Q
ec0f/g62676_db
ec0f/n_6701
ec0f/g62448_db
ec0f/n_3736
ec0f/g62512_sb
ec0f/g62676_sb
ec0f/g62676_da
ec0f/n_12337
ec0f/g64822_db
ec0f/g64822_da
ec0f/g62512_da
ec0f/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__37__Q
ec0f/n_7381
ec0f/g62512_db
ec0f/n_4905
ec0f/g64822_sb
ec0f/FE_OFN1440_n_12502
ec0f/n_1547
ec0f/n_12083
ec0f/n_11955
ec0f/n_7393
ec0f/n_5762
ec0f/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__2__Q
ec0f/n_6636
ec0f/g62476_sb
ec0f/n_11954
ec0f/FE_RN_425_0
ec0f/FE_RN_424_0
ec0f/g64839_db
ec0f/n_4441
ec0f/g62476_da
ec0f/g62476_db
ec0f/n_16445
ec0f/FE_OCP_RBN2009_FE_RN_290_0
ec0f/g67095_p
ec0f/n_11027
ec0f/n_12306
ec0f/n_6624
ec0f/n_10268
ec0f/n_16552
ec0f/n_16551
ec0f/g74944_p
ec0f/g64749_sb
ec0f/FE_OFN1792_n_4508
ec0f/n_10259
ec0f/n_16313
ec0f/FE_OFN1179_n_4143
ec0f/FE_OFN1180_n_4143
ec0f/FE_RN_290_0
ec0f/g74996_p
ec0f/n_15969
ec0f/n_16317
ec0f/g74943_p
ec0f/FE_RN_289_0
ec0f/FE_OCP_RBN2114_FE_RN_364_0
ec0f/n_9336
ec0f/FE_OFN964_n_4655
ec0f/g64915_db
ec0f/FE_OFN1428_n_12104
ec0f/n_10254
ec0f/n_12104
ec0f/n_9338
ec0f/g62613_db
ec0f/n_3688
ec0f/g64915_da
ec0f/g64915_sb
ec0f/n_4508
ec0f/n_10252
ec0f/g62613_sb
ec0f/g62613_da
ec0f/n_6331
ec0f/g62882_p
ec0f/FE_OFN1122_n_6935
ec0f/g66813_p
ec0f/FE_OFN1228_n_6624
ec0f/n_10780
ec0f/FE_OFN963_n_4655
ec0f/n_4655
ec0f/g67545_p
ec0f/n_6112
ec0f/n_1210
ec0f/n_4505
ec0f/n_1195
ec0f/g66658_p
ec0f/g66753_p
ec0f/n_4495
ec0f/FE_OFN623_n_4392
ec0f/n_4392
ec0f/n_1194
ec0f/n_4497
ec0f/n_242
ec0f/g67596_p
ec0f/g67493_p
ec0f/n_4409
ec0f/n_1106
ec0f/g66728_p
ec0f/n_1113
ec0f/g67390_p
ec0f/n_538
ec0f/n_4490
ec0f/g66627_p
ec0f/g64977_sb
ec0f/FE_OFN1456_n_12306
ec0f/g62392_db
ec0f/n_3594
ec0f/FE_OFN1730_n_11019
ec0f/g64977_da
ec0f/n_3650
ec0f/g64977_db
ec0f/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__6__Q
ec0f/g62392_sb
ec0f/g62392_da
ec0f/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__6__Q
ec0f/n_6814
ec0f/FE_OFN1528_n_4671
ec0f/g62516_db
ec0f/n_6546
ec0f/g62516_da
ec0f/g62516_sb
ec0f/g65099_da
ec0f/g65099_db
ec0f/n_11933
ec0f/g65099_sb
ec0f/g62675_db
ec0f/n_13310
ec0f/n_16589
ec0f/n_11932
ec0f/n_16588
ec0f/g64916_sb
ec0f/g64916_da
ec0f/g64974_sb
ec0f/FE_OFN1721_n_16317
ec0f/g62580_sb
ec0f/n_3687
ec0f/g64916_db
ec0f/n_6393
ec0f/g62580_da
ec0f/g62614_sb
ec0e/n_4306
ec0e/n_12321
ec0e/n_5916
ec0e/g62983_da
ec0e/g62983_sb
ec0e/g54346_sb
ec0e/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__11__Q
ec0e/n_5977
ec0e/g65417_sb
ec0e/g65417_da
ec0e/n_12753
ec0e/n_11842
ec0e/g64900_sb
ec0e/n_6238
ec0e/g62952_da
ec0e/g62952_db
ec0e/n_3512
ec0e/g65417_db
ec0e/g62586_db
ec0e/n_3693
ec0e/g64900_da
ec0e/g64900_db
ec0e/g62653_da
ec0e/g62952_sb
ec0e/n_6379
ec0e/g62586_da
ec0e/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__11__Q
ec0e/g62653_sb
ec0e/g65374_db
ec0e/n_11906
ec0e/n_12625
ec0e/n_12204
ec0e/g62586_sb
ec0e/n_12205
ec0e/g65374_sb
ec0e/g65374_da
ec0e/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__11__Q
ec0e/n_12876
ec0e/n_12626
ec0e/n_12875
ec0e/n_11905
ec0e/n_12488
ec0e/n_11904
ec0e/n_3529
ec0e/g62910_db
ec0e/n_6058
ec0e/g62337_sb
ec0e/g62337_da
ec0e/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__10__Q
ec0e/n_12624
ec0e/g62338_sb
ec0e/g62338_da
ec0e/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__11__Q
ec0e/g62910_da
ec0e/n_6924
ec0e/g62337_db
ec0e/n_3612
ec0e/n_6922
ec0e/g62338_db
ec0e/g62910_sb
ec0e/g64968_sb
ec0e/g65061_db
ec0e/n_12113
ec0e/n_3614
ec0e/g65059_db
ec0e/g64968_da
ec0e/g64968_db
ec0e/n_12755
ec0e/g65061_da
ec0e/g65061_sb
ec0e/n_12347
ec0e/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__11__Q
ec0e/g64861_db
ec0e/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__19__Q
ec0e/g64865_sb
ec0e/n_12437
ec0e/n_12416
ec0e/g62346_da
ec0e/g62346_sb
ec0e/g64861_da
ec0e/g64865_da
ec0e/n_4426
ec0e/g64865_db
ec0e/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__19__Q
ec0e/n_6908
ec0e/g62346_db
ec0e/n_4428
ec0e/g62688_db
ec0e/g62688_da
ec0e/g62688_sb
ec0e/g62522_da
ec0e/g62522_sb
ec0e/n_6657
ec0e/g62468_da
ec0e/g62468_sb
ec0e/n_6166
ec0e/g64858_db
ec0e/n_6532
ec0e/g62522_db
ec0e/g64858_sb
ec0e/g64858_da
ec0e/n_3718
ec0e/g62598_sb
ec0e/n_6900
ec0e/g62425_sb
ec0e/g62425_da
ec0e/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__27__Q
ec0e/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__21__Q
ec0e/n_6355
ec0e/g62598_da
ec0e/g62350_db
ec0e/n_3611
ec0e/g62350_da
ec0e/g62350_sb
ec0e/n_6747
ec0e/g62425_db
ec0e/n_4483
ec0e/g62598_db
ec0e/n_4325
ec0e/g65062_da
ec0e/g65062_db
ec0e/g62986_sb
ec0e/g64778_db
ec0e/g65046_da
ec0e/g65046_db
ec0e/g65062_sb
ec0e/g62986_da
ec0e/n_5910
ec0e/g64778_da
ec0e/g64778_sb
ec0e/g65046_sb
ec0e/g65333_db
ec0e/n_12305
ec0e/n_11838
ec0e/n_13314
ec0e/n_16600
ec0e/n_12275
ec0e/g64823_sb
ec0e/n_4264
ec0e/g65333_da
ec0e/n_17035
ec0e/n_12938
ec0e/n_17036
ec0e/g62916_sb
ec0e/n_13063
ec0e/FE_RN_380_0
ec0e/n_3735
ec0e/g64823_da
ec0e/g64823_db
ec0e/g65333_sb
ec0e/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__21__Q
ec0e/g63185_db
ec0e/g63185_sb
ec0e/n_12024
ec0e/n_12303
ec0e/FE_RN_379_0
ec0e/n_11990
ec0e/g62684_db
ec0e/n_5782
ec0e/g63185_da
ec0e/n_6171
ec0e/g62684_da
ec0e/g62684_sb
ec0e/g65362_db
ec0e/FE_OFN1724_n_14987
ec0e/g65301_db
ec0e/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__27__Q
ec0e/g63177_da
ec0e/g63177_sb
ec0e/FE_OFN1153_n_6391
ec0e/FE_OFN1158_n_6391
ec0e/n_3536
ec0e/g65362_da
ec0e/g63000_db
ec0e/n_5794
ec0e/g63177_db
ec0e/n_4275
ec0e/g65305_db
ec0e/g65362_sb
ec0e/g65305_da
ec0e/n_12660
ec0e/n_11941
ec0e/n_12895
ec0e/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__5__Q
ec0e/n_5985
ec0e/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__22__Q
ec0e/n_6580
ec0e/FE_OFN1178_n_4143
ec0e/g62501_da
ec0e/g62501_db
ec0e/g64782_da
ec0e/g64782_sb
ec0e/g62948_sb
ec0e/g62948_da
ec0e/g62948_db
ec0e/n_3532
ec0e/g62501_sb
ec0e/n_27
ec0e/n_3768
ec0e/g64782_db
ec0e/g65369_da
ec0e/g62359_db
ec0e/n_6880
ec0e/g62359_da
ec0g/n_13564
ec0g/wishbone_slave_unit_delayed_write_data_comp_wdata_out_92
ec0g/n_14316
ec0g/parchk_pci_ad_out_in_1190
ec0g/n_14377
ec0g/n_7661
ec0g/n_13290
ec0g/n_7307
ec0g/g53015_p
ec0g/n_13775
ec0g/n_13291
ec0g/n_13579
ec0g/FE_RN_136_0
ec0g/wishbone_slave_unit_delayed_write_data_comp_wdata_out_78
ec0g/g54231_db
ec0g/g54217_db
ec0g/n_13174
ec0g/g54217_da
ec0g/n_13572
ec0g/n_7502
ec0g/g53043_p
ec0g/n_13769
ec0g/FE_OFN1240_n_13668
ec0g/FE_OFN1661_n_13653
ec0g/g53931_db
ec0g/n_13162
ec0g/g54231_da
ec0g/g54140_da
ec0g/g54140_sb
ec0g/FE_OFN1666_n_13656
ec0g/n_13514
ec0g/g53931_da
ec0g/g54156_db
ec0g/wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_8__Q
ec0g/g53915_db
ec0g/g62064_sb
ec0g/g54156_sb
ec0g/n_7550
ec0g/FE_RN_135_0
ec0g/FE_OFN1665_n_13656
ec0g/n_14366
ec0g/n_7528
ec0g/n_13656
ec0g/g60339_p
ec0g/g53931_sb
ec0g/n_13237
ec0g/g54156_da
ec0g/g62064_da
ec0g/n_7745
ec0g/g62064_db
ec0g/g54244_da
ec0g/pci_target_unit_pci_target_if_pcir_fifo_ctrl_reg_77
ec0g/g54244_sb
ec0g/n_14374
ec0g/n_7655
ec0g/n_13443
ec0g/n_2123
ec0g/wishbone_slave_unit_pcim_sm_data_in_642
ec0g/n_13146
ec0g/parchk_pci_ad_out_in_1195
ec0g/g54140_db
ec0g/wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_22__Q
ec0g/g54131_db
ec0g/n_7637
ec0g/FE_OFN1662_n_13653
ec0g/g59722_p
ec0g/n_13527
ec0g/g53915_da
ec0g/n_13268
ec0g/n_14322
ec0g/n_14321
ec0g/g53915_sb
ec0g/g59345_p
ec0g/n_13765
ec0g/n_13569
ec0g/n_13571
ec0g/n_13347
ec0g/g62047_sb
ec0g/n_13578
ec0g/n_7548
ec0g/g53016_p
ec0g/n_13774
ec0g/n_13346
ec0g/g53087_p
ec0g/n_13768
ec0g/FE_RN_86_0
ec0g/FE_RN_84_0
ec0g/n_13460
ec0g/g62047_da
ec0g/n_14319
ec0g/g53098_p
ec0g/n_7636
ec0g/g62116_sb
ec0g/n_7764
ec0g/g62047_db
ec0g/wishbone_slave_unit_pcim_sm_data_in_656
ec0g/n_7553
ec0g/g53013_p
ec0g/n_14364
ec0g/n_14352
ec0g/n_2116
ec0g/g62119_sb
ec0g/parchk_pci_ad_out_in_1176
ec0g/n_14365
ec0g/n_7646
ec0g/n_7643
ec0g/FE_OFN923_n_13784
ec0g/n_13667
ec0g/g62115_sb
ec0g/g62115_da
ec0g/n_5579
ec0g/g62117_db
ec0g/n_17011
ec0g/FE_RN_365_0
ec0g/n_13289
ec0g/n_5581
ec0g/g62115_db
ec0g/FE_RN_366_0
ec0g/g53081_p
ec0g/n_13779
ec0g/FE_RN_367_0
ec0g/n_14373
ec0g/n_7654
ec0g/n_14320
ec0g/n_7634
ec0g/g53084_p
ec0g/n_14347
ec0g/n_7515
ec0g/parchk_pci_ad_out_in_1196
ec0g/FE_OFN1648_n_4868
ec0g/n_14348
ec0g/n_14376
ec0g/n_7660
ec0g/n_14378
ec0g/n_7663
ec0g/parchk_pci_ad_out_in_1189
ec0g/n_5585
ec0g/g62139_da
ec0g/g62139_sb
ec0g/g67100_p
ec0g/g67132_p
ec0g/g62112_db
ec0g/FE_OFN1649_n_4868
ec0g/n_14490
ec0g/parchk_pci_ad_out_in_1198
ec0g/n_5611
ec0g/g62094_da
ec0g/g62094_db
ec0g/g62094_sb
ec0g/n_667
ec0g/n_13831
ec0g/n_7658
ec0g/n_14531
ec0g/g66010_p
ec0g/n_605
ec0g/n_5554
ec0g/g62139_db
ec0g/g67102_p
ec0g/n_672
ec0g/g67145_p
ec0g/g67136_p
ec0g/n_1398
ec0g/g62099_da
ec0g/g62099_sb
ec0g/g62103_da
ec0g/g62103_sb
ec0g/g66004_p
ec0g/n_592
ec0g/g62093_da
ec0g/g62093_sb
ec0g/n_5604
ec0g/g62099_db
ec0g/n_5598
ec0g/g62103_db
ec0g/n_1403
ec0g/n_5612
ec0g/g62093_db
ec0g/g62100_sb
ec0g/g64381_p
ec0g/g62110_sb
ec0g/n_2252
ec0g/g64382_p
ec0g/n_1400
ec0g/g66008_p
ec0g/n_603
ec0h/n_2239
ec0h/n_1144
ec0h/pciu_bar1_in
ec0h/configuration_pci_err_data_512
ec0h/g67463_p
ec0h/n_7232
ec0h/n_6994
ec0h/n_14912
ec0h/n_7236
ec0h/n_15813
ec0h/n_2984
ec0h/g60614_db
ec0h/n_7429
ec0h/configuration_pci_err_data_509
ec0h/n_2836
ec0h/g67403_p
ec0h/n_1743
ec0h/n_7284
ec0h/pciu_am1_in_519
ec0h/FE_RN_409_0
ec0h/FE_RN_411_0
ec0h/FE_RN_410_0
ec0h/g66445_p
ec0h/n_439
ec0h/n_7484
ec0h/g60619_db
ec0h/g63268_p
ec0h/n_3406
ec0h/n_7483
ec0h/n_7055
ec0h/n_7453
ec0h/g67613_p
ec0h/n_7058
ec0h/n_5650
ec0h/n_3404
ec0h/n_4654
ec0h/pciu_bar1_in_381
ec0h/n_2927
ec0h/g60668_db
ec0h/n_5724
ec0h/n_2865
ec0h/n_15600
ec0h/n_15599
ec0h/n_4807
ec0h/n_4145
ec0h/FE_OCPN1989_n_16000
ec0h/n_3079
ec0h/n_3078
ec0h/FE_RN_400_0
ec0h/n_3070
ec0h/n_3292
ec0h/n_2821
ec0h/n_3042
ec0h/g65520_p
ec0h/n_2834
ec0h/n_2833
ec0h/n_6978
ec0h/n_4826
ec0h/n_3505
ec0h/FE_RN_401_0
ec0h/n_290
ec0h/n_5687
ec0h/g60642_db
ec0h/n_3403
ec0h/FE_OFN982_n_16720
ec0h/g61582_p
ec0h/n_4155
ec0h/g67495_p
ec0h/n_14919
ec0h/FE_RN_408_0
ec0h/FE_RN_406_0
ec0h/FE_RN_407_0
ec0h/g67505_p
ec0h/n_3039
ec0h/n_3288
ec0h/FE_OFN983_n_16720
ec0h/n_2857
ec0h/n_2856
ec0h/n_5643
ec0h/n_2621
ec0h/n_2840
ec0h/pciu_bar1_in_387
ec0h/n_17014
ec0h/g66449_p
ec0h/n_357
ec0h/pciu_am1_in_532
ec0h/pciu_bar1_in_394
ec0h/n_7494
ec0h/n_3232
ec0h/n_14934
ec0h/n_7049
ec0h/n_7477
ec0h/n_7439
ec0h/n_7068
ec0h/n_2076
ec0h/n_2830
ec0h/n_3424
ec0h/FE_OFN960_n_16810
ec0h/n_7486
ec0h/n_7059
ec0h/n_2074
ec0h/n_7255
ec0h/n_7254
ec0h/n_14926
ec0h/FE_OFN985_n_16720
ec0h/n_14929
ec0h/g63895_p
ec0h/n_7258
ec0h/n_7248
ec0h/n_2703
ec0h/n_2240
ec0h/FE_OFN961_n_16810
ec0h/n_3053
ec0h/n_2826
ec0h/n_7238
ec0h/n_7008
ec0h/n_7001
ec0h/FE_OCPN1974_FE_OFN961_n_16810
ec0h/n_7243
ec0h/n_3336
ec0h/n_1637
ec0h/n_4652
ec0h/n_6997
ec0h/n_2926
ec0h/n_3060
ec0h/n_2859
ec0h/n_6998
ec0h/n_3287
ec0h/n_3040
ec0h/n_2816
ec0h/g66441_p
ec0h/n_1148
ec0h/n_1141
ec0h/n_14925
ec0h/n_7251
ec0h/configuration_pci_err_data_523
ec0h/n_7285
ec0h/n_14931
ec0h/g66440_p
ec0h/n_302
ec0h/n_7458
ec0h/g66448_p
ec0h/n_436
ec0h/n_7002
ec0h/n_5669
ec0h/n_7229
ec0h/n_6993
ec0h/n_1149
ec0h/g67765_p
ec0h/pciu_bar1_in_393
ec0h/g60654_db
ec0h/n_4653
ec0h/n_3291
ec0h/n_3065
ec0h/n_7496
ec0h/pciu_bar0_in_370
ec0h/pciu_bar0_in_371
ec0h/n_3236
ec0h/g67783_p
ec0h/n_2913
ec0h/n_3062
ec0h/n_2775
ec0h/n_2082
ec0h/n_7069
ec0h/n_7579
ec0h/n_7407
ec0h/n_4808
ec0h/n_2843
ec0h/n_2802
ec0h/n_7404
ec0h/n_14928
ec0h/n_7576
ec0h/n_7414
ec0h/n_7585
ec0h/n_7246
ec0h/n_6999
ec0h/pciu_am1_in_535
ec0h/n_14927
ec0h/g67394_p
ec0h/n_7409
ec0h/pciu_am1_in_534
ec0h/n_225
ec0h/n_7581
ec0h/n_2286
ec0h/g67707_p
ec0h/pciu_bar1_in_397
ec0h/n_7247
ec0h/n_7000
ec0h/n_2077
ec0h/n_7413
ec0h/FE_OFN1001_n_7498
ec0h/n_7286
ec0h/n_7491
ec0h/n_7064
ec0h/n_1130
ec0h/n_7462
ec0h/n_7584
ec0h/n_7456
ec0h/g67329_p
ec0h/n_336
ec0h/g66451_p
ec0h/g66474_p
ec0h/n_227
ec0h/n_7245
ec0h/g67605_p
ec0h/g66442_p
ec0h/n_307
ec0h/n_7250
ec0h/n_7416
ec0h/n_431
ec0h/n_7435
ec0h/n_2083
ec0h/g67722_p
ec0h/n_7436
ec0h/n_7066
ech/n_15402
ech/FE_RN_14_0
ech/n_2883
ech/n_7319
ech/n_1617
ech/g59384_da
ech/FE_RN_240_0
ech/g66825_p
ech/parchk_pci_trdy_reg_in
ech/n_1618
ech/n_2370
ech/g59384_db
ech/wishbone_slave_unit_pcim_sm_last_in
ech/n_7539
ech/n_15799
ech/n_3081
ech/g64694_p
ech/n_2303
ech/g62319_p
ech/n_3450
ech/n_1192
ech/n_975
ech/n_2378
ech/n_4679
ech/g63307_p
ech/n_3023
ech/n_8532
ech/n_188
ech/n_3126
ech/n_7543
ech/n_1536
ech/n_6965
ech/n_1515
ech/pciu_pciif_stop_reg_in
ech/n_707
ech/wishbone_slave_unit_pci_initiator_sm_timeout
ech/n_3127
ech/n_8752
ech/n_8749
ech/n_8750
ech/n_378
ech/wishbone_slave_unit_pci_initiator_sm_transfer
ech/n_2132
ech/wbu_pciif_frame_out_in
ech/n_3378
ech/g65555_p
ech/n_1514
ech/pci_target_unit_pcit_if_comp_flush_in
ech/FE_OFN740_n_2746
ech/n_3812
ech/n_2726
ech/n_2043
ech/n_3163
ech/g65493_p
ech/g64707_p
ech/n_3379
ech/n_16496
ech/n_2803
ech/n_2443
ech/n_1964
ech/g66854_p
ech/pci_target_unit_del_sync_comp_flush_out_reg_Q
ech/n_1459
ech/wishbone_slave_unit_pci_initiator_sm_mabort2
ech/n_2805
ech/n_4792
ech/n_7210
ech/configuration_meta_cache_lsize_to_wb_bits_929
ech/n_2951
ech/n_3408
ech/n_2900
ech/n_3260
ech/n_4793
ech/pciu_cache_line_size_in_776
ech/n_3047
ech/n_15406
ech/n_1615
ech/g74154_p
ech/n_7400
ech/configuration_meta_cache_lsize_to_wb_bits_927
ech/configuration_sync_cache_lsize_to_wb_bits_reg_4__Q
ech/n_1616
ech/FE_RN_20_0
ech/pci_target_unit_pci_target_sm_rd_from_fifo
ech/g67369_p
ech/pciu_cache_line_size_in_777
ech/pciu_cache_line_size_in_775
ech/FE_RN_19_0
ech/FE_RN_18_0
ech/FE_RN_12_0
ech/n_15401
ech/n_532
ech/configuration_meta_cache_lsize_to_wb_bits_928
ech/FE_OFN739_n_2746
ech/n_2747
ech/FE_RN_13_0
ech/n_1126
ech/n_15400
ech/g67745_p
ech/FE_OFN178_n_7210
ech/n_2746
ech/pci_target_unit_pci_target_if_target_rd_completed
ech/n_2287
ech/n_1088
ech/n_2887
ech/FE_OCPN1848_n_16798
ech/n_2374
ech/g65995_db
ech/n_2046
ech/n_3380
ech/FE_OFN1104_n_7400
ech/pci_target_unit_pci_target_sm_state_transfere_reg
ech/n_1450
ech/n_152
ech/n_2765
ech/FE_OFN1483_n_15366
ech/pci_target_unit_pci_target_sm_state_transfere_reg_reg_Q
ech/FE_RN_225_0
ech/n_2147
ech/g66001_da
ech/g66001_db
ech/FE_OFN192_n_2683
ech/n_205
ech/n_2718
ech/g66000_da
ech/g66000_db
ech/g67082_db
ech/n_454
ech/FE_OFN188_n_1193
ech/g60697_sb
ech/g67082_da
ech/n_47
ech/n_2683
ech/n_1505
ech/g67092_db
ech/n_1193
ech/g60697_da
ech/g67082_sb
ech/parchk_pci_irdy_en_in
ech/n_447
ech/out_bckp_irdy_out
ech/n_2471
ech/g60697_db
ech/n_2946
ech/n_16330
ech/FE_RN_28_0
ech/n_16328
ech/FE_RN_29_0
ech/n_8539
ech/parchk_pci_frame_en_in
ech/FE_RN_27_0
ech/n_16329
ech/g74961_p
ech/n_15366
ech/g74434_db
ech/n_8574
ech/n_2351
ech/pci_target_unit_pci_target_sm_previous_frame
ech/g65996_db
ech/n_2372
ech/g74434_da
ech/FE_OFN1482_n_15366
ech/g74434_sb
h0a/n_896
h0a/n_1373
h0a/n_897
h0a/n_1974
h0a/n_1374
h0a/n_977
h0a/g66138_p
h0a/n_1986
h0a/n_1987
h0a/n_1985
h0a/n_2930
h0a/n_1975
h0a/n_1477
h0a/g65261_p
h0a/n_2224
h0a/n_563
h0a/n_562
h0a/g67519_p
h0a/pci_target_unit_fifos_pciw_addr_data_in_124
h0a/n_16292
h0a/n_16304
h0a/n_14856
h0a/n_14858
h0a/n_14770
h0a/g64597_p
h0a/g65523_p
h0a/n_13377
h0a/n_14863
h0a/n_14780
h0a/n_14708
h0a/n_14642
h0a/pci_target_unit_fifos_pciw_addr_data_in_129
h0a/n_14577
h0a/n_208
h0a/pci_target_unit_fifos_pciw_addr_data_in_144
h0a/n_14625
h0a/n_14668
h0a/n_14761
h0a/n_14849
h0a/n_13367
h0a/n_15196
h0a/n_15197
h0a/n_15187
h0a/n_14730
h0a/n_14658
h0a/n_16231
h0a/n_3873
h0a/g64302_da
h0a/g64302_db
h0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__5__Q
h0a/g64302_sb
h0a/g63085_da
h0a/g63085_sb
h0a/n_5084
h0a/g63085_db
h0a/FE_OFN1021_g64577_p
h0a/n_16240
h0a/n_14635
h0a/n_14699
h0a/n_14580
h0a/n_14409
h0a/n_14499
h0a/FE_OFN1020_g64577_p
h0a/g64347_sb
h0a/g64347_da
h0a/n_3830
h0a/g63013_sb
h0a/g64347_db
h0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__9__Q
h0a/n_5076
h0a/g63089_db
h0a/g63089_da
h0a/g63089_sb
h0a/n_3869
h0a/g64306_da
h0a/g64306_db
h0a/g64306_sb
h0a/n_13923
h0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__9__Q
h0a/g63052_db
h0a/n_5146
h0a/g63052_da
h0a/g64265_da
h0a/g64265_sb
h0a/n_3908
h0a/g63052_sb
h0a/g64265_db
h0a/n_16261
h0a/g62773_sb
h0a/g62773_db
h0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__9__Q
h0a/g62773_da
h0a/n_4001
h0a/n_5448
h0a/g64164_db
h0a/g64164_da
h0a/g64164_sb
h0a/g64261_sb
h0a/g64261_db
h0a/n_3912
h0a/g64261_da
h0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__5__Q
h0a/g63047_da
h0a/g63047_sb
h0a/n_5158
h0a/g63047_db
h0a/n_13930
h0a/g64120_sb
h0a/g64120_da
h0a/g62853_sb
h0a/n_4040
h0a/g64120_db
h0a/g62853_da
h0a/g53297_p
h0a/n_13849
h0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__5__Q
h0a/g62853_db
h0a/n_5263
h0a/g53298_p
h0a/g62833_sb
h0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__11__Q
h0a/n_5308
h0a/g62833_da
h0a/n_4005
h0a/g64160_db
h0a/g62833_db
h0a/g64160_da
h0a/g64160_sb
h0a/g64197_sb
h0a/g64197_da
h0a/g62843_sb
h0a/n_3972
h0a/g64197_db
h0a/g62843_da
h0a/g62843_db
h0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__11__Q
h0a/n_5285
h0a/n_13846
h0a/g53313_p
h0a/n_14400
h0a/n_16616
h0a/n_16617
h0a/g53314_p
h0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__9__Q
h0a/n_5283
h0a/g62844_db
h0a/g62844_da
h0a/g64199_db
h0a/n_3970
h0a/g62844_sb
h0a/g64199_da
h0a/g64199_sb
h0a/g64253_db
h0a/n_17022
h0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__9__Q
h0a/g64253_sb
h0a/g64253_da
h0a/n_3920
h0a/g63096_da
h0a/g63096_sb
h0a/g63096_db
h0a/n_5062
h0a/g63165_sb
h0a/g64366_db
h0a/g63165_da
h0a/n_3814
h0a/g64366_da
h0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__5__Q
h0a/g64366_sb
h0a/n_14097
h0a/n_5476
h0a/g62752_da
h0a/g62752_db
h0a/g64105_db
h0a/n_13904
h0a/n_14298
h0a/n_14067
h0a/n_14477
h0a/n_14243
h0a/n_14245
h0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__11__Q
h0a/g64083_db
h0a/g62811_db
h0a/n_5356
h0a/g62811_da
h0a/g62720_db
h0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__9__Q
h0a/n_5543
h0a/g62720_da
h0a/g64205_db
h0a/n_14165
h0a/n_14164
h0a/g64205_sb
h0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__9__Q
h0a/n_5511
h0a/g62734_da
h0a/g62734_db
h0a/n_14016
h0a/n_14401
h0a/n_13863
h0a/n_14493
h0a/g64352_db
h0a/g64352_sb
h0a/n_17023
h0a/g64352_da
h0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__9__Q
h0a/n_4965
h0a/g63141_da
h0a/n_3826
h0a/g63141_sb
h0a/g63141_db
h0a/g64129_da
h0a/g64129_sb
h0a/FE_OFN1056_g64577_p
h0a/g64129_db
h0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__7__Q
h0a/n_4033
h0a/g62851_da
h0a/g62851_sb
h0a/n_4957
h0a/g63165_db
h0a/n_14592
h0a/FE_OFN1576_n_16657
h0a/g62752_sb
h0a/n_4052
h0a/g64105_da
h0a/g64105_sb
h0a/g64157_sb
h0a/g64307_da
h0a/g64307_sb
h0a/g64307_db
h0a/g64206_da
h0a/g64206_sb
h0a/g64083_da
h0a/g64083_sb
h0a/n_4072
h0a/g62811_sb
h0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__7__Q
h0a/n_5523
h0a/g62728_db
h0a/g62728_da
h0a/g62728_sb
h0a/n_4026
h0a/g62720_sb
h0a/n_3964
h0a/g64136_db
h0a/g64205_da
h0a/g64136_da
h0a/g64136_sb
h0a/FE_OFN1039_g64577_p
h0a/FE_OFN1049_g64577_p
h0a/FE_OCPN1924_FE_OFN1758_n_13997
h0a/FE_OCP_RBN2088_FE_OFN1756_n_13997
h0a/g62734_sb
h0a/n_4044
h0a/g64116_da
h0a/g64116_db
h0a/g64116_sb
h0a/FE_OFN971_n_4727
h0a/g64093_sb
h0a/g64093_da
h0a/n_16257
h0a/n_14018
h0a/n_13865
h0a/n_4062
h0a/g64093_db
h0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__7__Q
h0a/g62810_da
h0a/g62810_sb
h0a/g62810_db
h0a/n_5358
h0a/n_5267
h0a/g62851_db
h0a/g64085_da
h0a/g64085_sb
h0a/n_4070
h0a/g64085_db
h0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__4__Q
h0a/g62759_da
h0a/g62759_sb
h0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__11__Q
h0a/n_5265
h0a/g62818_sb
h0a/g62852_db
h0a/g62852_da
h0a/g64221_da
h0a/g64221_sb
h0a/g64206_db
h0a/n_3963
h0a/g62852_sb
h0a/g64134_da
h0a/g64134_sb
h0a/n_14597
h0a/FE_OFN1769_n_13800
h0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__7__Q
h0a/n_5269
h0a/g62850_da
h0a/g62850_db
h0a/n_14169
h0a/n_14168
h0a/g74886_p
h0a/n_16255
h0a/n_16260
h0a/n_16258
h0a/n_4968
h0a/g63140_da
h0a/g63140_db
h0a/g64361_sb
h0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__7__Q
h0a/g64361_da
h0a/n_13926
h0a/n_16256
h0a/n_13925
h0a/g64321_sb
h0a/g64321_da
h0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__7__Q
h0a/g63143_db
h0a/n_4961
h0a/g63143_da
h0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__4__Q
h0a/n_5205
h0a/g63021_db
h0a/g63021_da
h0a/g64236_da
h0a/g64236_sb
h0a/n_3936
h0a/g64236_db
h0a/g63021_sb
h0a/n_14173
h0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__4__Q
h0a/FE_OFN1775_n_13971
h0a/g62759_db
h0a/n_5472
h0a/n_14174
h0a/g64119_sb
h0a/g62818_db
h0a/g62818_da
h0a/n_3948
h0a/n_5339
h0a/g64221_db
h0a/g64134_db
h0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__26__Q
h0a/n_4028
h0a/n_5429
h0a/g62781_da
h0a/g62781_db
h0a/g62781_sb
h0a/n_5080
h0a/g63087_da
h0a/g63087_db
h0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__7__Q
h0a/g63087_sb
h0a/g62850_sb
h0a/n_3871
h0a/n_3966
h0a/g64203_da
h0a/g64203_db
h0a/g64304_da
h0a/g64304_db
h0a/g64304_sb
h0a/g64203_sb
h0a/FE_OFN1014_g64577_p
h0a/n_16259
h0a/g63049_sb
h0a/g63049_da
h0a/n_3910
h0a/g63049_db
h0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__7__Q
h0a/g64361_db
h0a/g63140_sb
h0a/n_3818
h0a/g64263_da
h0a/g64263_sb
h0a/g64263_db
h0a/FE_OCP_RBN2079_n_16975
h0a/g64321_db
h0a/n_3855
h0a/g63143_sb
h0a/n_5086
h0a/g63084_da
h0a/g63084_db
h0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__4__Q
h0a/n_14100
h0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__4__Q
h0a/n_13931
h0a/FE_OFN1025_g64577_p
h0a/g64098_sb
h0a/g64098_da
h0a/n_16232
h0a/n_14099
h0a/n_16238
h0a/n_13932
h0a/n_16234
h0a/n_16239
h0a/n_16237
h0a/n_16233
h0a/g63046_sb
h0a/g62824_db
h0a/g63046_da
h0a/n_3913
h0a/g64092_sb
h0a/g64092_da
h0a/g64260_db
h0a/g64260_da
h0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__4__Q
h0a/g64260_sb
h0a/n_5330
h0a/g62824_da
h0a/FE_OFN1551_n_4732
h0a/n_4063
h0a/g64092_db
h0a/g64350_sb
h0a/g64350_da
h0a/g64350_db
h0a/n_3828
h0a/g63070_da
h0a/g63070_sb
h0a/FE_OFN1045_g64577_p
h0a/n_5110
h0a/g63070_db
h0a/g64100_sb
h0a/g64100_da
h0a/n_4055
h0a/g64100_db
h0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__19__Q
h0a/g62815_da
h0a/g62815_sb
h0a/n_13927
h0a/n_13928
h0a/n_5153
h0a/g64341_db
h0a/g64317_sb
h0a/g64317_db
h0a/g64341_sb
h0a/g64317_da
h0a/n_3859
h0a/g63084_sb
h0a/n_4947
h0a/g63176_db
h0a/g63176_da
h0a/g64098_db
h0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__4__Q
h0a/n_4057
h0a/g62741_da
h0a/g62741_sb
h0a/n_5497
h0a/g62741_db
h0a/g63046_db
h0a/n_5161
h0a/g64159_sb
h0a/g64159_da
h0a/FE_OFN1606_n_4740
h0a/g64279_db
h0a/g63062_sb
h0a/n_3894
h0a/g64279_da
h0a/g63062_da
h0a/FE_OFN1031_g64577_p
h0a/g64279_sb
h0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__19__Q
h0a/n_13982
h0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__19__Q
h0a/n_5126
h0a/g63062_db
h0a/n_13981
h0a/n_16220
h0a/n_14226
h0a/n_14055
h0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__19__Q
h0a/n_5347
h0a/g62815_db
h0a/n_5235
h0a/FE_OFN972_n_4727
h0a/g63028_sb
h0a/g63028_da
h0a/n_3837
h0a/g64285_db
h0a/g64341_da
h0a/g64285_sb
h0a/FE_OFN947_n_4725
h0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__24__Q
h0a/n_5190
h0a/g63028_db
h0a/n_13970
h0a/g64357_sb
h0a/g64357_da
h0a/g63176_sb
h0a/n_3821
h0a/g64357_db
h0a/FE_OFN1605_n_4740
h0a/n_14022
h0a/n_16236
h0a/n_16235
h0a/n_13868
h0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__4__Q
h0a/g64144_db
h0a/g62823_da
h0a/n_4020
h0a/g62823_sb
h0a/g64144_da
h0a/g64144_sb
h0a/g62812_sb
h0a/g62812_da
h0a/n_4006
h0a/g64159_db
h0a/n_5354
h0a/g62812_db
h0a/n_3946
h0a/g64223_db
h0a/g64240_db
h0a/n_3932
h0a/g64240_da
h0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__19__Q
h0a/g63023_sb
h0a/g64240_sb
h0a/g63023_da
h0a/n_5298
h0a/g62838_da
h0a/g62838_db
h0a/n_5200
h0a/g63023_db
h0a/n_16223
h0a/n_16222
h0a/n_16221
h0a/g64180_sb
h0a/g64180_da
h0a/g64180_db
h0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__19__Q
h0a/n_3986
h0a/g64167_sb
h0a/g64167_da
h0a/g62790_da
h0a/g62790_sb
h0a/n_3998
h0a/g64167_db
h0a/n_5409
h0a/g62790_db
h0a/g62865_da
h0a/g62865_sb
h0a/g62865_db
h0a/g64334_db
h0a/g63068_sb
h0a/n_3888
h0a/g64285_da
h0a/g63068_da
h0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__24__Q
h0a/n_5114
h0a/g63068_db
h0a/n_13969
h0a/n_16229
h0a/n_16230
h0a/n_16228
h0a/n_16227
h0a/g74859_p
h0a/FE_OFN1577_n_16657
h0a/n_14044
h0a/n_13887
h0a/FE_OFN948_n_4725
h0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__24__Q
h0a/FE_OCP_RBN2078_n_16975
h0a/n_5404
h0a/g62792_db
h0a/g62792_da
h0a/g62823_db
h0a/n_5332
h0a/g64118_da
h0a/g64118_sb
h0a/g64118_db
h0a/n_4042
h0a/g64162_sb
h0a/g62838_sb
h0a/g64258_sb
h0a/g64258_db
h0a/n_3915
h0a/g64258_da
h0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__19__Q
h0a/g63102_da
h0a/g63102_sb
h0a/n_14142
h0a/n_14960
h0a/n_14961
h0a/n_14144
h0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__19__Q
h0a/g64254_db
h0a/n_3919
h0a/g64254_da
h0a/g64254_sb
h0a/g63038_da
h0a/g63038_sb
h0a/g63131_sb
h0a/g63131_da
h0a/n_3843
h0a/n_4988
h0a/g63131_db
h0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__24__Q
h0a/g64334_da
h0a/g64334_sb
h0a/g63107_sb
h0a/g63107_db
h0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__24__Q
h0a/g63107_da
h0a/n_3861
h0a/n_5040
h0a/g64314_da
h0a/g64314_db
h0a/g64314_sb
h0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__24__Q
h0a/n_5258
h0a/g62855_db
h0a/g62855_da
h0a/g64137_db
h0a/n_4025
h0a/g62855_sb
h0a/g64137_da
h0a/g64137_sb
h0a/g62792_sb
h0a/g64292_da
h0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__31__Q
h0a/g64292_sb
h0a/n_3881
h0a/g64292_db
h0a/FE_OFN1036_g64577_p
h0a/n_5050
h0a/g63102_db
h0a/g64198_da
h0a/g64198_sb
h0a/n_3971
h0a/g64198_db
h0a/g62841_sb
h0a/g62841_da
h0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__20__Q
h0a/n_5290
h0a/g62841_db
h0a/g63038_db
h0a/n_5172
h0a/g64287_db
h0a/FE_OFN1030_g64577_p
h0a/g64161_db
h0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__27__Q
h0a/g64161_sb
h0a/g64161_da
h0a/n_4004
h0a/n_5337
h0a/g62819_da
h0a/g62819_db
h0a/g62819_sb
h0a/n_14130
h0a/n_16225
h0a/n_14129
h0a/g64173_da
h0a/g64173_sb
h0a/n_16226
h0a/g63037_sb
h0a/g63037_da
h0a/n_3840
h0a/g64337_da
h0a/g64337_db
h0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__31__Q
h0a/g64337_sb
h0a/n_13956
h0a/g53250_p
h0a/n_13853
h0a/n_14250
h0a/n_5098
h0a/g63076_da
h0a/g63076_db
h0a/g62766_db
h0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__31__Q
h0a/g63076_sb
h0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__27__Q
h0a/n_5240
h0a/g62863_da
h0a/g62863_db
h0a/g62863_sb
h0a/n_3951
h0a/n_14203
h0a/g64218_db
h0a/g64218_da
h0a/n_14205
h0a/n_14447
h0a/g64218_sb
h0a/g64089_da
h0a/g64089_sb
h0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__27__Q
h0a/n_5108
h0a/n_16625
h0a/n_14260
h0a/g63071_db
h0a/n_13965
h0a/n_13963
h0a/g63071_da
h0a/n_16624
h0a/n_14446
h0a/n_3886
h0a/g63071_sb
h0a/g64287_da
h0a/g64287_sb
h0a/g53230_p
h0a/g53231_p
h0a/n_13884
h0a/n_14041
h0a/g63111_db
h0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__27__Q
h0a/n_5033
h0a/g63111_da
h0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__27__Q
h0a/n_3858
h0a/g63111_sb
h0a/n_5433
h0a/g64318_da
h0a/g64318_sb
h0a/g62779_db
h0a/g64318_db
h0a/g62779_da
h0a/g64173_db
h0a/n_3992
h0a/g62779_sb
h0a/g64087_da
h0a/g64087_sb
h0a/n_14212
h0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__24__Q
h0a/n_14211
h0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__24__Q
h0a/n_5174
h0a/g63037_db
h0a/g64088_db
h0a/n_4067
h0a/g64088_da
h0a/g64088_sb
h0a/n_14435
h0a/g53251_p
h0a/n_14034
h0a/n_13879
h0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__31__Q
h0a/n_5463
h0a/g64250_db
h0a/g64250_sb
h0a/g64250_da
h0a/n_4034
h0a/g62771_sb
h0a/g64128_db
h0a/g64128_da
h0a/g64128_sb
h0a/g64089_db
h0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__20__Q
h0a/g62816_da
h0a/n_4066
h0a/g62816_sb
h0a/pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__27__Q
h0a/n_5183
h0a/g63032_db
h0a/g63032_da
h0a/g64342_sb
h0a/g64248_da
h0a/g64248_sb
h0a/g63032_sb
h0a/n_3924
h0a/g64248_db
h0a/n_14124
h0a/n_14123
h0a/g64335_da
h0a/g64335_sb
h0a/n_3842
h0a/g64335_db
h0a/g62730_sb
h0a/g62730_da
h0a/n_4068
h0a/g64087_db
h0a/n_5519
h0a/g62730_db
h0a/n_5499
h0a/g62740_db
h0a/g62740_da
h0a/g62740_sb
h0a/g64086_da
h0a/g64086_sb
h0a/n_5396
h0a/g62795_db
h0a/g62795_da
h0a/g64181_db
h0a/n_3985
h0a/g62795_sb
h0a/g64181_da
h0a/g64181_sb
h0a/g63026_da
h0a/g63026_sb
h0a/n_5194
h0a/g63026_db
h0a/n_5345
h0a/g62816_db
h0a/g64342_db
h0a/n_3836
h0a/g64342_da
h0a/g63024_sb
h0a/g63133_sb
h0a/g64228_db
h0a/g64228_sb
h0a/g64228_da
h0a/n_5470
h0a/g62762_db
h0a/g62762_da
h0a/g64086_db
h0a/n_4069
h0a/g62764_da
h0a/g62764_sb
h0a/n_5467
h0a/g62764_db
h0b/g62418_da
h0b/g62418_sb
h0b/FE_OCP_RBN2075_n_11767
h0b/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__17__Q
h0b/n_6301
h0b/g62627_da
h0b/g62627_db
h0b/g62627_sb
h0b/g62462_da
h0b/g62462_sb
h0b/n_6672
h0b/g62462_db
h0b/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__13__Q
h0b/n_6680
h0b/FE_RN_54_0
h0b/g62588_db
h0b/n_4411
h0b/g64901_db
h0b/n_4410
h0b/g64901_da
h0b/g64901_sb
h0b/FE_OFN1439_n_12502
h0b/g64840_sb
h0b/n_6761
h0b/g62418_db
h0b/g64978_db
h0b/n_4367
h0b/g64978_da
h0b/g64978_sb
h0b/g64924_sb
h0b/g64924_da
h0b/n_4391
h0b/g64924_db
h0b/g62459_sb
h0b/g64830_db
h0b/n_4451
h0b/g64830_da
h0b/g64830_sb
h0b/g64828_sb
h0b/g64828_da
h0b/g64828_db
h0b/n_4453
h0b/g62458_db
h0b/g62458_da
h0b/g62458_sb
h0b/FE_RN_56_0
h0b/FE_RN_55_0
h0b/n_12780
h0b/g62588_sb
h0b/n_6374
h0b/g62588_da
h0b/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__13__Q
h0b/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__247
h0b/n_12448
h0b/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__13__Q
h0b/g65405_db
h0b/g65405_sb
h0b/g65405_da
h0b/n_3518
h0b/n_12654
h0b/n_12361
h0b/n_5928
h0b/g62977_sb
h0b/g62977_da
h0b/g62977_db
h0b/g63144_sb
h0b/n_4239
h0b/g65396_da
h0b/g65396_sb
h0b/g65396_db
h0b/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__14__Q
h0b/n_6308
h0b/g62624_sb
h0b/g62624_da
h0b/g62624_db
h0b/g65073_db
h0b/n_4309
h0b/g65073_da
h0b/g65073_sb
h0b/g62459_da
h0b/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__14__Q
h0b/n_6678
h0b/g62459_db
h0b/g65071_db
h0b/n_4311
h0b/g65071_da
h0b/g65071_sb
h0b/g62548_sb
h0b/g62548_db
h0b/n_3657
h0b/n_6470
h0b/g62548_da
h0b/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__6__Q
h0b/g64961_da
h0b/g64961_db
h0b/g64961_sb
h0b/g62369_db
h0b/n_4492
h0b/n_6865
h0b/g62369_da
h0b/g62369_sb
h0b/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__0__Q
h0b/g62584_sb
h0b/g62584_db
h0b/n_4368
h0b/g64975_da
h0b/g64975_db
h0b/g62584_da
h0b/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__0__Q
h0b/n_6384
h0b/n_12519
h0b/n_12003
h0b/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__24__Q
h0b/g63144_da
h0b/n_5852
h0b/g63144_db
h0b/g65355_da
h0b/g65355_sb
h0b/n_4317
h0b/g65355_db
h0b/g64995_sb
h0b/g64995_db
h0b/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__0__Q
h0b/g64995_da
h0b/n_4356
h0b/n_6806
h0b/g62397_da
h0b/g62397_sb
h0b/g62397_db
h0b/n_12339
h0b/g62401_sb
h0b/FE_OFN1735_n_12004
h0b/g62401_da
h0b/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__13__Q
h0b/n_6797
h0b/g62401_db
h0b/n_4321
h0b/n_12063
h0b/g65052_da
h0b/g65052_db
h0b/g65052_sb
h0b/g64804_sb
h0b/g64804_da
h0b/g62382_sb
h0b/g62382_db
h0b/n_4463
h0b/g64804_db
h0b/n_6837
h0b/g62382_da
h0b/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__24__Q
h0b/n_12869
h0b/g62651_sb
h0b/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__0__Q
h0b/n_6243
h0b/g62651_da
h0b/g62651_db
h0b/n_4360
h0b/g64761_sb
h0b/g64761_da
h0b/g64761_db
h0b/g64988_da
h0b/g64988_db
h0b/g64988_sb
h0b/n_11913
h0b/n_11912
h0b/FE_RN_375_0
h0b/n_12286
h0b/g64975_sb
h0b/n_12810
h0b/n_11914
h0b/n_11915
h0b/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__0__Q
h0b/g65347_da
h0b/g65347_sb
h0b/g63147_da
h0b/g63147_sb
h0b/n_5846
h0b/g63147_db
h0b/n_4259
h0b/g65401_db
h0b/g65401_sb
h0b/g65401_da
h0b/FE_OFN1526_n_4671
h0b/n_11916
h0b/n_12213
h0b/g65344_sb
h0b/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__0__Q
h0b/g65344_db
h0b/g65344_da
h0b/n_4261
h0b/n_6031
h0b/g62925_da
h0b/g62925_sb
h0b/g62925_db
h0b/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__13__Q
h0b/n_6311
h0b/g62623_da
h0b/g62623_db
h0b/FE_RN_385_0
h0b/FE_RN_387_0
h0b/FE_RN_386_0
h0b/FE_RN_390_0
h0b/g64922_db
h0b/n_4393
h0b/g64922_da
h0b/g64922_sb
h0b/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__9__Q
h0b/n_6323
h0b/g62617_sb
h0b/g62617_da
h0b/g62617_db
h0b/n_3636
h0b/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__243
h0b/n_3637
h0b/g65010_db
h0b/g65010_da
h0b/g65010_sb
h0b/g62667_sb
h0b/g62667_db
h0b/n_4342
h0b/g62667_da
h0b/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__24__Q
h0b/n_6204
h0b/g65017_db
h0b/n_12284
h0b/n_12720
h0b/g62990_sb
h0b/n_13064
h0b/n_12927
h0b/g65347_db
h0b/g62680_sb
h0b/g65051_db
h0b/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__6__Q
h0b/g62680_db
h0b/n_3619
h0b/g65051_da
h0b/g65051_sb
h0b/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__0__Q
h0b/n_5856
h0b/g63094_da
h0b/g63094_db
h0b/g63094_sb
h0b/n_4247
h0b/g65378_da
h0b/g65378_sb
h0b/g65378_db
h0b/FE_RN_389_0
h0b/FE_RN_388_0
h0b/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__13__Q
h0b/g65407_sb
h0b/g65407_da
h0b/n_4232
h0b/g65407_db
h0b/g62623_sb
h0b/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__13__Q
h0b/g65366_sb
h0b/g65366_da
h0b/n_4252
h0b/g65366_db
h0b/FE_RN_376_0
h0b/n_12460
h0b/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__260
h0b/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__26__Q
h0b/n_6345
h0b/n_4403
h0b/g62603_da
h0b/g62603_db
h0b/n_4404
h0b/g64909_db
h0b/g62603_sb
h0b/g64909_da
h0b/n_12450
h0b/g62999_sb
h0b/g62999_da
h0b/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__4__Q
h0b/g65017_sb
h0b/g65017_da
h0b/g62999_db
h0b/n_4253
h0b/n_5884
h0b/FE_RN_374_0
h0b/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__26__Q
h0b/n_5902
h0b/g62990_da
h0b/g62990_db
h0b/g65384_da
h0b/g65384_sb
h0b/n_4656
h0b/g65384_db
h0b/g62680_da
h0b/g65363_db
h0b/n_6179
h0b/g63002_db
h0b/n_3535
h0b/g65363_da
h0b/g65363_sb
h0b/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__7__Q
h0b/n_12212
h0b/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_13_
h0b/n_4280
h0b/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__0__Q
h0b/n_6061
h0b/g65294_db
h0b/n_5816
h0b/g63160_sb
h0b/g63160_da
h0b/g63160_db
h0b/g62433_sb
h0b/g62928_sb
h0b/g62928_da
h0b/n_6025
h0b/g62928_db
h0b/g64914_da
h0b/g64914_sb
h0b/n_4397
h0b/g64914_db
h0b/g62612_db
h0b/n_4396
h0b/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__238
h0b/g64909_sb
h0b/n_12452
h0b/n_12785
h0b/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__9__Q
h0b/g65361_da
h0b/g65361_sb
h0b/g63004_sb
h0b/g65361_db
h0b/g63004_da
h0b/n_5874
h0b/g63004_db
h0b/n_3534
h0b/g65365_da
h0b/g65365_sb
h0b/g65365_db
h0b/n_5878
h0b/g63002_da
h0b/g63002_sb
h0b/g62962_sb
h0b/g62962_db
h0b/n_4224
h0b/g62908_sb
h0b/g65294_sb
h0b/g62908_da
h0b/g65424_db
h0b/g65294_da
h0b/g62908_db
h0b/n_4281
h0b/n_4236
h0b/g65402_da
h0b/g65402_db
h0b/g62939_db
h0b/g62939_sb
h0b/n_12610
h0b/n_11801
h0b/n_12611
h0b/n_12340
h0b/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__14__Q
h0b/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__14__Q
h0b/g62894_da
h0b/g62894_sb
h0b/g62433_da
h0b/n_6731
h0b/g62433_db
h0b/g64812_db
h0b/n_4461
h0b/g65379_db
h0b/n_4246
h0b/g65379_da
h0b/g64812_da
h0b/g65379_sb
h0b/g62968_db
h0b/g64812_sb
h0b/n_6333
h0b/g62612_da
h0b/g62612_sb
h0b/n_5946
h0b/g62968_da
h0b/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__4__Q
h0b/g62968_sb
h0b/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__4__Q
h0b/g65308_db
h0b/n_4272
h0b/g65308_da
h0b/g62922_db
h0b/n_6037
h0b/g62922_da
h0b/g62922_sb
h0b/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__4__Q
h0b/g65308_sb
h0b/g63161_sb
h0b/g63161_db
h0b/n_3569
h0b/g65311_db
h0b/g65311_da
h0b/g65311_sb
h0b/g63161_da
h0b/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__7__Q
h0b/n_5814
h0b/g65312_db
h0b/g65312_sb
h0b/g65312_da
h0b/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__9__Q
h0b/n_3568
h0b/g63154_db
h0b/n_5833
h0b/g63154_da
h0b/g62962_da
h0b/n_6647
h0b/g62472_da
h0b/g62472_sb
h0b/g65424_da
h0b/g65424_sb
h0b/n_13049
h0b/g65402_sb
h0b/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__26__Q
h0b/n_6003
h0b/g62939_da
h0b/n_12279
h0b/g65278_sb
h0b/g65278_da
h0b/g62894_db
h0b/n_4288
h0b/n_6089
h0b/g65278_db
h0b/g54596_p
h0b/g65074_sb
h0b/g65074_da
h0b/n_3605
h0b/g65074_db
h0b/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__25__Q
h0b/g62442_db
h0b/n_11944
h0b/g62551_sb
h0b/g62551_db
h0b/n_3658
h0b/g62551_da
h0b/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__9__Q
h0b/n_6463
h0b/n_11942
h0b/n_12498
h0b/g62970_sb
h0b/g65343_db
h0b/g62970_db
h0b/n_3545
h0b/g65343_da
h0b/g62970_da
h0b/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__9__Q
h0b/g65343_sb
h0b/n_5942
h0b/n_11918
h0b/n_12882
h0b/n_12636
h0b/n_12490
h0b/n_11919
h0b/n_12637
h0b/n_12353
h0b/n_12219
h0b/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__8__Q
h0b/n_5868
h0b/g63007_da
h0b/g63007_sb
h0b/g63007_db
h0b/n_4267
h0b/g65326_da
h0b/g65326_sb
h0b/g65326_db
h0b/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__14__Q
h0b/n_6795
h0b/g62402_sb
h0b/g62402_da
h0b/g62402_db
h0b/g64789_db
h0b/n_4477
h0b/g64789_da
h0b/g64789_sb
h0b/g64837_sb
h0b/g64837_da
h0b/n_12400
h0b/n_6712
h0b/g62442_da
h0b/g62442_sb
h0b/g64960_sb
h0b/g64960_da
h0b/g62682_db
h0b/n_4324
h0b/g64960_db
h0b/g65048_da
h0b/g65048_db
h0b/n_4323
h0b/g65048_sb
h0b/n_12812
h0b/n_12499
h0b/g64785_sb
h0b/g64785_da
h0b/n_3766
h0b/g64785_db
h0b/g62710_db
h0b/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__9__Q
h0b/n_6150
h0b/g62710_da
h0b/g62710_sb
h0b/n_11924
h0b/g65075_sb
h0b/g65075_da
h0b/n_3604
h0b/g65075_db
h0b/g62400_db
h0b/n_13051
h0b/n_12712
h0b/n_11995
h0b/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__26__Q
h0b/g62927_sb
h0b/n_6929
h0b/g62335_sb
h0b/g62335_da
h0b/g62335_db
h0b/g62927_db
h0b/n_4194
h0b/g64795_db
h0b/g65314_db
h0b/n_4469
h0b/g64795_da
h0b/g64795_sb
h0b/g65004_sb
h0b/g65004_da
h0b/g54591_p
h0b/g64837_db
h0b/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__25__Q
h0b/n_3728
h0b/n_12094
h0b/n_6649
h0b/g62471_db
h0b/g62471_da
h0b/g62471_sb
h0b/g65089_sb
h0b/g65089_da
h0b/g54594_p
h0b/g62682_sb
h0b/g65089_db
h0b/g62682_da
h0b/n_6175
h0b/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__359
h0b/g62394_da
h0b/g62394_sb
h0b/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__8__Q
h0b/n_6184
h0b/g62678_da
h0b/g62678_db
h0b/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__4__Q
h0b/g62678_sb
h0b/g64757_db
h0b/n_11946
h0b/g64783_sb
h0b/g64783_da
h0b/n_3767
h0b/g64783_db
h0b/g62400_da
h0b/g62400_sb
h0b/g62927_da
h0b/n_3639
h0b/n_4301
h0b/g62394_db
h0b/n_4499
h0b/g64757_da
h0b/g64757_sb
h1a/n_12202
h1a/n_12208
h1a/g65321_db
h1a/g65367_db
h1a/n_4416
h1a/g64884_db
h1a/n_12201
h1a/n_12623
h1a/n_3567
h1a/n_12874
h1a/g65313_da
h1a/g65313_sb
h1a/g65313_db
h1a/g62455_sb
h1a/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__10__Q
h1a/n_6686
h1a/g62455_da
h1a/g62553_sb
h1a/g62553_da
h1a/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__10__Q
h1a/n_6458
h1a/g62553_db
h1a/n_12348
h1a/n_13309
h1a/n_13048
h1a/n_3708
h1a/g64879_da
h1a/g64879_db
h1a/g64879_sb
h1a/g62697_sb
h1a/g62697_da
h1a/n_6160
h1a/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__11__Q
h1a/n_6607
h1a/g62489_sb
h1a/g62489_da
h1a/g62489_db
h1a/n_3633
h1a/n_15439
h1a/n_12207
h1a/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__30__Q
h1a/n_5995
h1a/g62943_da
h1a/g62943_db
h1a/n_3561
h1a/g65321_da
h1a/g65321_sb
h1a/g62943_sb
h1a/g65367_sb
h1a/g65367_da
h1a/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__18__Q
h1a/n_6017
h1a/n_4251
h1a/g62932_da
h1a/g62932_sb
h1a/g62932_db
h1a/n_16407
h1a/n_13067
h1a/g54569_p
h1a/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__18__Q
h1a/n_6440
h1a/g62560_da
h1a/g62560_db
h1a/g62560_sb
h1a/n_16403
h1a/n_16406
h1a/n_16402
h1a/g62561_sb
h1a/g62561_da
h1a/n_6438
h1a/g62561_db
h1a/n_16404
h1a/n_11841
h1a/n_5966
h1a/n_12752
h1a/g65298_db
h1a/n_3575
h1a/g65298_da
h1a/g63167_db
h1a/g62958_da
h1a/g62958_db
h1a/g62958_sb
h1a/g63167_sb
h1a/n_5804
h1a/g63167_da
h1a/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__16__Q
h1a/g65315_sb
h1a/g65315_db
h1a/g65315_da
h1a/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__16__Q
h1a/n_3566
h1a/n_6021
h1a/g62930_da
h1a/g62930_db
h1a/g62930_sb
h1a/n_12783
h1a/n_12463
h1a/n_12877
h1a/n_12206
h1a/n_11908
h1a/n_11806
h1a/n_12349
h1a/n_11903
h1a/n_11805
h1a/n_12203
h1a/n_12345
h1a/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__10__Q
h1a/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__10__Q
h1a/n_6610
h1a/g65018_db
h1a/g62488_sb
h1a/g62488_da
h1a/g62488_db
h1a/g65018_da
h1a/g65018_sb
h1a/g54586_p
h1a/g64843_db
h1a/n_3726
h1a/g64843_da
h1a/g64843_sb
h1a/n_13317
h1a/n_13068
h1a/n_12253
h1a/g54568_p
h1a/n_12759
h1a/n_12326
h1a/n_12325
h1a/n_12044
h1a/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_12__487
h1a/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__19__Q
h1a/n_28
h1a/n_6789
h1a/n_12528
h1a/n_4472
h1a/g64792_da
h1a/g64792_db
h1a/g64792_sb
h1a/n_12943
h1a/n_12047
h1a/n_12751
h1a/n_12750
h1a/n_11971
h1a/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__18__Q
h1a/n_6592
h1a/n_12318
h1a/n_12045
h1a/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__19__Q
h1a/n_6589
h1a/g62916_db
h1a/g62497_sb
h1a/g62497_da
h1a/g65008_db
h1a/g62497_db
h1a/n_6047
h1a/n_4349
h1a/g65008_da
h1a/g65008_sb
h1a/g65298_sb
h1a/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__16__Q
h1a/n_5824
h1a/n_11888
h1a/n_12182
h1a/n_12598
h1a/g65087_sb
h1a/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__16__Q
h1a/g54606_p
h1a/n_12859
h1a/n_12480
h1a/n_11885
h1a/n_13042
h1a/n_16401
h1a/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__10__Q
h1a/n_6318
h1a/g62620_da
h1a/g62620_db
h1a/g65076_db
h1a/g62620_sb
h1a/n_6315
h1a/g62621_da
h1a/g62621_db
h1a/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__11__Q
h1a/g62621_sb
h1a/g64810_sb
h1a/g64810_da
h1a/g64810_db
h1a/n_3748
h1a/g62429_db
h1a/n_12908
h1a/n_12682
h1a/n_11972
h1a/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__30__Q
h1a/n_12684
h1a/n_12683
h1a/n_12946
h1a/g62405_sb
h1a/g62405_da
h1a/g62405_db
h1a/g64831_sb
h1a/g64831_da
h1a/n_12758
h1a/n_12757
h1a/g64832_sb
h1a/n_12323
h1a/n_12252
h1a/g62496_sb
h1a/g62496_da
h1a/g62496_db
h1a/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__30__Q
h1a/n_4435
h1a/g64848_db
h1a/g64848_da
h1a/g64848_sb
h1a/g65301_sb
h1a/g63157_db
h1a/n_3554
h1a/g63157_da
h1a/g64963_sb
h1a/g63157_sb
h1a/g65330_da
h1a/g65330_db
h1a/g65330_sb
h1a/n_16399
h1a/n_12935
h1a/n_12059
h1a/n_12058
h1a/n_12596
h1a/n_12335
h1a/n_12481
h1a/n_11798
h1a/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__16__Q
h1a/n_6087
h1a/g62895_da
h1a/g62895_db
h1a/g62895_sb
h1a/n_3603
h1a/g65076_da
h1a/g65076_sb
h1a/g63162_sb
h1a/g63162_da
h1a/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__10__Q
h1a/g64918_sb
h1a/g64918_da
h1a/n_3685
h1a/g64918_db
h1a/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__11__Q
h1a/n_6741
h1a/n_6093
h1a/g62892_da
h1a/g62892_sb
h1a/g62892_db
h1a/g62429_da
h1a/g62429_sb
h1a/g64970_sb
h1a/g64970_da
h1a/n_3653
h1a/g64970_db
h1a/g62417_db
h1a/n_6763
h1a/g62417_da
h1a/g62417_sb
h1a/g62463_sb
h1a/n_6670
h1a/g62463_da
h1a/g62463_db
h1a/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__18__Q
h1a/n_4449
h1a/g64831_db
h1a/n_12108
h1a/n_12418
h1a/g64832_da
h1a/g64832_db
h1a/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__19__Q
h1a/n_4448
h1a/n_12107
h1a/g62464_db
h1a/n_12415
h1a/n_6668
h1a/g62464_da
h1a/g62464_sb
h1a/g62510_sb
h1a/g62510_da
h1a/n_6558
h1a/g62510_db
h1a/g64990_db
h1a/n_3646
h1a/g64990_da
h1a/n_16400
h1a/n_16398
h1a/g64963_da
h1a/n_3656
h1a/g64963_db
h1a/g62343_db
h1a/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__16__Q
h1a/n_6913
h1a/g62343_da
h1a/g62343_sb
h1a/n_12421
h1a/n_12597
h1a/g64956_sb
h1a/g64956_da
h1a/g65279_sb
h1a/g65279_da
h1a/n_3585
h1a/g65279_db
h1a/g65368_db
h1a/n_5812
h1a/g63162_db
h1a/n_3587
h1a/g65276_da
h1a/g65276_sb
h1a/g65276_db
h1a/g65410_sb
h1a/g65410_da
h1a/n_3640
h1a/g65410_db
h1a/n_3516
h1a/g65001_da
h1a/g65001_db
h1a/g65001_sb
h1a/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__30__Q
h1a/g65287_da
h1a/g65287_sb
h1a/n_3581
h1a/g65287_db
h1a/n_5792
h1a/g63178_db
h1a/g63178_da
h1a/g63178_sb
h1a/g65273_sb
h1a/g62897_sb
h1a/g65273_da
h1a/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__19__Q
h1a/g62897_da
h1a/g62897_db
h1a/n_4291
h1a/g65273_db
h1a/n_6083
h1a/g64926_sb
h1a/g64926_da
h1a/g64926_db
h1a/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__19__Q
h1a/g64953_sb
h1a/g64953_da
h1a/g64953_db
h1a/n_4377
h1a/g62437_db
h1a/n_6722
h1a/g62437_da
h1a/g62437_sb
h1a/n_16397
h1a/g64990_sb
h1a/g62665_db
h1a/n_3668
h1a/n_6208
h1a/g62665_da
h1a/g62665_sb
h1a/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__22__Q
h1a/g64948_db
h1a/n_12299
h1a/n_12735
h1a/g64956_db
h1b/g65859_db
h1b/g61948_sb
h1b/g61948_da
h1b/n_1580
h1b/g65859_da
h1b/g65676_da
h1b/g65676_sb
h1b/g65815_db
h1b/FE_OFN905_n_2055
h1b/g65815_sb
h1b/n_1901
h1b/g65815_da
h1b/pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__23__Q
h1b/g61867_sb
h1b/g61867_da
h1b/g65676_db
h1b/n_7929
h1b/g61948_db
h1b/pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__3__Q
h1b/g65859_sb
h1b/n_8102
h1b/g61867_db
h1b/g62005_sb
h1b/g65965_db
h1b/g62005_da
h1b/n_2158
h1b/g65965_da
h1b/n_7885
h1b/g62005_db
h1b/g65965_sb
h1b/pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__23__Q
h1b/n_11091
h1b/n_11093
h1b/n_11092
h1b/g61813_db
h1b/pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__23__Q
h1b/n_8166
h1b/g61813_da
h1b/pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__23__Q
h1b/g61813_sb
h1b/g65798_db
h1b/n_1665
h1b/g65818_db
h1b/g61871_sb
h1b/n_1898
h1b/g65818_da
h1b/g61871_da
h1b/g65798_da
h1b/g65818_sb
h1b/pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__27__Q
h1b/g65758_db
h1b/g65798_sb
h1b/n_2045
h1b/g65758_da
h1b/g65758_sb
h1b/g65966_db
h1b/g62009_sb
h1b/n_16585
h1b/pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__27__Q
h1b/g62009_db
h1b/g61871_db
h1b/n_8092
h1b/n_2157
h1b/g65966_da
h1b/g62009_da
h1b/n_7877
h1b/g65966_sb
h1b/g65949_db
h1b/g65836_db
h1b/g65949_sb
h1b/n_1562
h1b/g65949_da
h1b/pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__23__Q
h1b/pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__23__Q
h1b/n_1883
h1b/g65836_da
h1b/g65836_sb
h1b/g61902_sb
h1b/g61902_da
h1b/g61936_da
h1b/g61936_sb
h1b/n_8019
h1b/g61902_db
h1b/g65710_db
h1b/pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__7__Q
h1b/n_7951
h1b/g61936_db
h1b/g65710_da
h1b/g65710_sb
h1b/g65771_sb
h1b/g65845_db
h1b/g65771_da
h1b/g65789_db
h1b/pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__7__Q
h1b/n_1875
h1b/g65845_da
h1b/g65845_sb
h1b/g61917_sb
h1b/n_1602
h1b/g65771_db
h1b/pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__7__Q
h1b/g61828_sb
h1b/g61917_da
h1b/g61828_da
h1b/pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__7__Q
h1b/g65789_sb
h1b/g62020_sb
h1b/g62020_da
h1b/n_2152
h1b/g65972_db
h1b/g65972_da
h1b/n_7855
h1b/g62020_db
h1b/pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__7__Q
h1b/g65972_sb
h1b/g61917_db
h1b/g61828_db
h1b/n_7987
h1b/n_8130
h1b/n_10781
h1b/pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__7__Q
h1b/n_11043
h1b/pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__7__Q
h1b/n_8208
h1b/g65722_db
h1b/n_8064
h1b/g65881_da
h1b/g65881_sb
h1b/g61883_db
h1b/g61795_db
h1b/g61795_da
h1b/g65722_sb
h1b/g61883_da
h1b/g65722_da
h1b/n_1940
h1b/n_1865
h1b/g65881_db
h1b/g61883_sb
h1b/g61795_sb
h1b/g65739_sb
h1b/n_11780
h1b/pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__31__Q
h1b/n_7999
h1b/g61911_da
h1b/g61911_db
h1b/g65842_da
h1b/g65842_sb
h1b/g61911_sb
h1b/n_1878
h1b/g65842_db
h1b/g61946_db
h1b/n_7933
h1b/g65773_sb
h1b/g65773_da
h1b/g65773_db
h1b/n_1912
h1b/g61758_da
h1b/g61758_sb
h1b/FE_OFN1061_n_8407
h1b/n_1957
h1b/g61791_sb
h1b/g61791_da
h1b/n_8218
h1b/g61791_db
h1b/n_8246
h1b/g61780_db
h1b/g61780_da
h1b/g61780_sb
h1b/n_8288
h1b/g61762_sb
h1b/g61762_db
h1b/g61762_da
h1b/n_1945
h1b/n_11774
h1b/n_8362
h1b/g61729_db
h1b/g61729_da
h1b/n_2189
h1b/g61729_sb
h1b/g65789_da
h1b/g65862_db
h1b/g65862_sb
h1b/g65862_da
h1b/pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__7__Q
h1b/n_11042
h1b/n_1707
h1b/g61952_da
h1b/g61952_sb
h1b/n_7921
h1b/g61952_db
h1b/g65739_db
h1b/pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__31__Q
h1b/g61789_db
h1b/n_8223
h1b/g61789_da
h1b/n_1932
h1b/g65739_da
h1b/g61789_sb
h1b/g62014_sb
h1b/g62014_db
h1b/g62014_da
h1b/g65914_db
h1b/n_8297
h1b/g61758_db
h1b/g65735_sb
h1b/g65735_da
h1b/g65708_sb
h1b/g65708_da
h1b/n_1947
h1b/g65708_db
h1b/g61784_sb
h1b/g61784_da
h1b/pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__27__Q
h1b/n_8236
h1b/g61784_db
h1b/pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__31__Q
h1b/n_8302
h1b/g61756_sb
h1b/g61756_db
h1b/g61756_da
h1b/n_2039
h1b/g65683_db
h1b/n_11778
h1b/pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__31__Q
h1b/g65683_da
h1b/g65695_db
h1b/n_2205
h1b/g65695_da
h1b/g65683_sb
h1b/g65695_sb
h1b/g65786_sb
h1b/g65786_da
h1b/g65786_db
h1b/pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__31__Q
h1b/n_1598
h1b/g61822_sb
h1b/g61822_da
h1b/n_8144
h1b/g61822_db
h1b/n_11063
h1b/n_11064
h1b/g65742_sb
h1b/FE_OFN1060_n_8407
h1b/g65821_db
h1b/g65821_sb
h1b/n_1895
h1b/g65821_da
h1b/g61876_da
h1b/g61876_sb
h1b/g61876_db
h1b/g61940_sb
h1b/n_1568
h1b/g65914_da
h1b/pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__27__Q
h1b/g65914_sb
h1b/g61940_da
h1b/g61940_db
h1b/n_7943
h1b/n_1608
h1b/g65735_db
h1b/g61817_sb
h1b/g61817_da
h1b/g65839_db
h1b/pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__27__Q
h1b/n_1880
h1b/g65839_da
h1b/pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__27__Q
h1b/g65839_sb
h1b/n_8157
h1b/g61817_db
h1b/n_11079
h1b/n_16586
h1b/g65751_sb
h1b/g65751_da
h1b/g65707_da
h1b/g65707_sb
h1b/n_2061
h1b/g65707_db
h1b/pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__27__Q
h1b/g61718_db
h1b/n_8389
h1b/g61718_da
h1b/g61718_sb
h1b/g61723_db
h1b/n_8376
h1b/n_1571
h1b/g65900_da
h1b/g65900_db
h1b/g61723_da
h1b/pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__28__Q
h1b/g65900_sb
h1b/g61723_sb
h1b/g65887_sb
h1b/g65887_da
h1b/pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__28__Q
h1b/g61907_da
h1b/n_1862
h1b/g61907_sb
h1b/g65887_db
h1b/pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__30__Q
h1b/n_8226
h1b/g61788_db
h1b/g61788_da
h1b/g65742_db
h1b/n_1929
h1b/g61788_sb
h1b/g65742_da
h1b/g61821_db
h1b/pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__30__Q
h1b/g61821_sb
h1b/g65820_db
h1b/g65820_sb
h1b/n_1896
h1b/g65820_da
h1b/g61875_sb
h1b/g65823_sb
h1b/n_1893
h1b/g65823_da
h1b/pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__6__Q
h1b/g61882_da
h1b/g61882_sb
h1b/n_8066
h1b/g61882_db
h1b/g61906_sb
h1b/g61906_da
h1b/n_8009
h1b/g61906_db
h1b/n_1923
h1b/g65751_db
h1b/g61751_sb
h1b/n_11081
h1b/g61751_da
h1b/pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__27__Q
h1b/n_8313
h1b/g61751_db
h1b/g61941_sb
h1b/g61941_da
h1b/n_7941
h1b/g61941_db
h1b/n_11076
h1b/g61907_db
h1b/n_8007
h1b/g65804_db
h1b/pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__28__Q
h1b/n_1906
h1b/g65804_da
h1b/g65804_sb
h1b/g61785_da
h1b/g61785_sb
h1b/n_10782
h1b/g65698_sb
h1b/n_8147
h1b/g65698_da
h1b/g61821_da
h1b/g65806_db
h1b/n_1589
h1b/g65806_da
h1b/g65806_sb
h1b/n_11067
h1b/g62019_da
h1b/g62019_sb
h1b/g62019_db
h1b/n_7857
h1b/g65851_db
h1b/n_2184
h1b/g65851_da
h1b/g65851_sb
h1b/pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__10__Q
h1b/g61991_sb
h1b/g61991_da
h1b/n_7913
h1b/g61991_db
h1b/g62025_sb
h1b/g65750_sb
h1b/g65750_da
h1b/n_1605
h1b/g65750_db
h1b/g61799_da
h1b/g61799_sb
h1b/g65797_sb
h1b/g65797_da
h1b/g61818_sb
h1b/n_1591
h1b/g65797_db
h1b/g61818_da
h1b/g65747_sb
h1b/pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__28__Q
h1b/n_8154
h1b/g61818_db
h1b/n_11075
h1b/n_8234
h1b/g61785_db
h1b/g65953_sb
h1b/g65953_da
h1b/pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__28__Q
h1b/g65953_db
h1b/n_2167
h1b/g62010_da
h1b/g62010_sb
h1b/g65698_db
h1b/pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__30__Q
h1b/n_2203
h1b/g61722_sb
h1b/g61722_da
h1b/g61819_sb
h1b/n_8379
h1b/g61722_db
h1b/g65874_db
h1b/g65874_da
h1b/pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__9__Q
h1b/g65874_sb
h1b/n_1869
h1b/g61919_db
h1b/g61919_da
h1b/g61919_sb
h1b/pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__10__Q
h1b/n_7847
h1b/g65868_sb
h1b/g65868_da
h1b/g62025_da
h1b/g62025_db
h1b/n_2054
h1b/g65868_db
h1b/n_11153
h1b/pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__10__Q
h1b/n_8198
h1b/g61799_db
h1b/g65731_sb
h1b/g65731_da
h1b/pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__28__Q
h1b/n_8311
h1b/g65747_da
h1b/g61752_da
h1b/g61752_db
h1b/n_1925
h1b/g61752_sb
h1b/g65747_db
h1b/n_11078
h1b/n_11077
h1b/g65706_sb
h1b/n_2200
h1b/g65706_da
h1b/g65706_db
h1b/g61719_da
h1b/g61719_sb
h1b/pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__28__Q
h1b/g65908_db
h1b/n_1855
h1b/g65908_da
h1b/g65908_sb
h1b/n_7875
h1b/g62010_db
h1b/g61819_db
h1b/pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__29__Q
h1b/n_8152
h1b/g61819_da
h1b/n_1604
h1b/g65755_da
h1b/g65755_db
h1b/g65755_sb
h1b/g65906_db
h1b/g65906_da
h1b/g65906_sb
h1b/FE_OFN915_n_2053
h1b/n_7983
h1b/pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__10__Q
h1b/n_8054
h1b/FE_RN_320_0
h1b/FE_RN_322_0
h1b/FE_RN_321_0
h1b/pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__10__Q
h1b/n_8279
h1b/g61766_db
h1b/g61766_da
h1b/g65731_db
h1b/g65775_sb
h1b/g65775_da
h1b/n_1936
h1b/g61766_sb
h1b/n_2192
h1b/g65775_db
h1b/g61700_sb
h1b/g61700_da
h1b/pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__10__Q
h1b/n_8428
h1b/g61700_db
h1b/pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__28__Q
h1b/g61719_db
h1b/n_8387
h1b/n_8089
h1b/g61872_db
h1b/g61872_da
h1b/g61872_sb
h1b/g65935_db
h1b/n_2169
h1b/g65935_da
h1b/g62012_da
h1b/g62012_sb
h1b/g65682_sb
h1b/g65682_da
h1b/pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__29__Q
h1b/g65682_db
h1b/n_1955
h1b/g61786_da
h1b/g61786_sb
h1b/n_8231
h1b/g61786_db
h1b/g61830_db
h1b/n_8125
h1b/g65848_sb
h1b/g65848_da
h1b/pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__10__Q
h1b/n_7979
h1b/n_1587
h1b/g65848_db
h1b/g61921_da
h1b/g61921_db
h1b/g61921_sb
h1b/n_11147
h1b/n_11796
h1b/n_11155
h1b/g65690_da
h1b/g65690_sb
h1b/n_1953
h1b/g65690_db
h1b/g61733_sb
h1b/g65854_sb
h1b/g61944_db
h1b/g61944_da
h1b/g65854_da
h1b/n_1702
h1b/g61944_sb
h1b/g65854_db
h1b/g65841_sb
h1b/g65841_da
h1b/n_8003
h1b/g61909_db
h1b/g61909_da
h1b/g65841_db
h1b/n_1879
h1b/g61909_sb
h1b/g65935_sb
h1b/g62012_db
h1b/n_7871
h1b/g65738_sb
h1b/n_2056
h1b/g65738_da
h1b/g65738_db
h1b/g61793_sb
h1c/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__7__Q
h1c/n_6065
h1c/g62906_db
h1c/n_3578
h1c/n_11812
h1c/g65419_da
h1c/g65419_sb
h1c/n_4227
h1c/g65419_db
h1c/g62453_db
h1c/n_3733
h1c/g65082_db
h1c/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__0__Q
h1c/n_6743
h1c/g62428_da
h1c/g62428_sb
h1c/g62619_da
h1c/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__0__Q
h1c/g62906_da
h1c/g65290_da
h1c/g65290_sb
h1c/g62483_sb
h1c/g62483_da
h1c/n_6321
h1c/g62619_db
h1c/n_4302
h1c/g65088_db
h1c/g63155_db
h1c/n_4270
h1c/g65088_da
h1c/g65320_sb
h1c/n_12489
h1c/n_12068
h1c/g65324_da
h1c/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__6__Q
h1c/g65324_sb
h1c/g65290_db
h1c/g65088_sb
h1c/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_2__6
h1c/FE_RN_295_0
h1c/FE_RN_296_0
h1c/g64825_sb
h1c/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__6__Q
h1c/g64825_db
h1c/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__9__Q
h1c/g64825_da
h1c/n_12072
h1c/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__7__Q
h1c/n_6691
h1c/g62453_da
h1c/g62453_sb
h1c/g62648_sb
h1c/n_6252
h1c/g64939_db
h1c/g62648_db
h1c/n_3675
h1c/g62481_sb
h1c/n_4338
h1c/g64964_sb
h1c/g65320_da
h1c/g65320_db
h1c/g63155_sb
h1c/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__24__Q
h1c/n_3559
h1c/g65324_db
h1c/g64840_db
h1c/g62648_da
h1c/g62449_sb
h1c/g62449_db
h1c/n_4375
h1c/g64964_da
h1c/g64964_db
h1c/g62947_da
h1c/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__4__Q
h1c/g62947_sb
h1c/FE_OFN1749_n_11027
h1c/n_5830
h1c/g63155_da
h1c/n_5827
h1c/g63156_db
h1c/n_12635
h1c/n_3734
h1c/g64824_da
h1c/g64824_db
h1c/g64824_sb
h1c/g62451_sb
h1c/g62530_db
h1c/n_3758
h1c/n_6514
h1c/g62530_sb
h1c/n_6398
h1c/g62578_da
h1c/g62578_db
h1c/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__4__Q
h1c/g62578_sb
h1c/n_4359
h1c/n_6699
h1c/g62449_da
h1c/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__4__Q
h1c/n_5987
h1c/g62947_db
h1c/n_4519
h1c/g65370_da
h1c/g65370_sb
h1c/g65370_db
h1c/g63156_sb
h1c/g63156_da
h1c/n_12005
h1c/n_12352
h1c/n_12067
h1c/g62530_da
h1c/g64798_db
h1c/n_11947
h1c/g64989_db
h1c/n_12076
h1c/n_12402
h1c/n_12366
h1c/n_12664
h1c/n_12666
h1c/n_11948
h1c/n_12235
h1c/g62454_db
h1c/n_4455
h1c/g62454_da
h1c/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__0__Q
h1c/g62454_sb
h1c/g65021_sb
h1c/n_6689
h1c/g62486_db
h1c/n_3632
h1c/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__7__Q
h1c/g64798_da
h1c/g65325_sb
h1c/n_12521
h1c/n_12006
h1c/g64798_sb
h1c/n_12663
h1c/g62707_sb
h1c/g64826_db
h1c/g62451_db
h1c/n_6695
h1c/g62451_da
h1c/g65021_da
h1c/g62949_sb
h1c/n_12724
h0c/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__17__Q
h0c/n_6911
h0c/g62543_da
h0c/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__31__Q
h0c/g62543_sb
h0c/n_5872
h0c/g63005_da
h0c/g63005_db
h0c/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__36__Q
h0c/g63005_sb
h0c/g62344_da
h0c/n_4394
h0c/g62344_sb
h0c/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__1__Q
h0c/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__56
h0c/n_12479
h0c/n_6480
h0c/g62344_db
h0c/g64815_da
h0c/g64815_sb
h0c/g64815_db
h0c/g64920_da
h0c/g64920_sb
h0c/n_4395
h0c/g64920_db
h0c/n_12475
h0c/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__70
h0c/n_12809
h0c/g62361_sb
h0c/g64873_da
h0c/g64873_sb
h0c/n_12792
h0c/g65921_da
h0c/g65921_sb
h0c/n_1850
h0c/g64801_da
h0c/g64801_db
h0c/g64801_sb
h0c/n_4422
h0c/g64873_db
h0c/g62543_db
h0c/g65921_db
h0c/n_12378
h0c/n_2379
h0c/g65671_da
h0c/g65671_db
h0c/g65671_sb
h0c/g62438_da
h0c/g62438_sb
h0c/FE_OFN1155_n_6391
h0c/n_6720
h0c/g62438_db
h0c/n_3743
h0c/n_4313
h0c/g65068_da
h0c/g65068_db
h0c/n_4312
h0c/g62478_db
h0c/n_4333
h0c/g65034_sb
h0c/n_6631
h0c/g62478_da
h0c/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__31__Q
h0c/g62478_sb
h0c/n_6127
h0c/g62755_da
h0c/g62755_db
h0c/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__36__Q
h0c/g62755_sb
h0c/g62945_da
h0c/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__36__Q
h0c/g62945_sb
h0c/n_11957
h0c/n_11956
h0c/g65057_sb
h0c/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__31__Q
h0c/n_6876
h0c/g65068_sb
h0c/g62361_da
h0c/g62361_db
h0c/g65034_da
h0c/g65034_db
h0c/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__17__Q
h0c/n_6724
h0c/g62436_sb
h0c/g62436_da
h0c/g62436_db
h0c/n_4319
h0c/g65057_da
h0c/g65057_db
h0c/g62711_da
h0c/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__31__Q
h0c/g62711_sb
h0c/n_6148
h0c/n_12419
h0c/g62711_db
h0c/n_4307
h0c/g65080_da
h0c/g65080_db
h0c/n_12080
h0c/n_12679
h0c/n_12380
h0c/g62945_db
h0c/n_1852
h0c/n_5991
h0c/g65916_da
h0c/g65916_sb
h0c/g65916_db
h0c/n_4456
h0c/g64820_da
h0c/g64820_db
h0c/g64820_sb
h0c/n_11981
h0c/g62432_sb
h0c/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__13__Q
h0c/n_6733
h0c/g62432_da
h0c/g62432_db
h0c/n_4316
h0c/g65063_da
h0c/g65063_db
h0c/g65063_sb
h0c/n_12766
h0c/n_12110
h0c/n_12343
h0c/n_12949
h0c/n_12964
h0c/n_12950
h0c/n_12767
h0c/g62896_db
h0c/n_4289
h0c/g65275_da
h0c/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__17__Q
h0c/g65275_sb
h0c/g65080_sb
h0c/g65275_db
h0c/g64935_da
h0c/g64935_sb
h0c/FE_OFN1172_n_4093
h0c/n_4384
h0c/g64935_db
h0c/n_6144
h0c/g62713_da
h0c/g62713_sb
h0c/g62713_db
h0c/n_5864
h0c/g63009_db
h0c/n_6053
h0c/g62913_da
h0c/g62913_db
h0c/g62913_sb
h0c/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__17__Q
h0c/n_5969
h0c/g62956_da
h0c/g62956_db
h0c/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__17__Q
h0c/n_4221
h0c/g62956_sb
h0c/n_12051
h0c/n_6085
h0c/g62896_da
h0c/g62896_sb
h0c/n_5993
h0c/g62944_da
h0c/g62944_db
h0c/n_12618
h0c/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__31__Q
h0c/g62944_sb
h0c/n_12906
h0c/n_13055
h0c/n_12505
h0c/n_4269
h0c/g65322_da
h0c/g65322_db
h0c/g62642_db
h0c/n_6264
h0c/g62642_da
h0c/n_11980
h0c/g62642_sb
h0c/n_11892
h0c/g65329_db
h0c/n_4266
h0c/g65329_da
h0c/n_5772
h0c/g63192_da
h0c/g63192_db
h0c/g65400_da
h0c/g65400_sb
h0c/n_4237
h0c/g65400_db
h0c/n_4220
h0c/g65434_da
h0c/g65434_db
h0c/g65433_da
h0c/g65433_sb
h0c/g65434_sb
h0c/g65433_db
h0c/n_12331
h0c/g62524_da
h0c/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__13__Q
h0c/g62524_sb
h0c/n_11843
h0c/n_12764
h0c/g62524_db
h0c/n_4370
h0c/g65036_da
h0c/g65036_sb
h0c/n_4332
h0c/g65036_db
h0c/g62340_sb
h0c/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__13__Q
h0c/g62340_db
h0c/n_6919
h0c/g62340_da
h0c/n_11969
h0c/g65322_sb
h0c/g62508_da
h0c/g62508_sb
h0c/n_6563
h0c/g62508_db
h0c/n_16596
h0c/g63184_da
h0c/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__13__Q
h0c/g63192_sb
h0c/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__13__Q
h0c/n_5973
h0c/g62954_db
h0c/n_4249
h0c/g62954_da
h0c/g62954_sb
h0c/g65375_da
h0c/g65375_db
h0c/g65375_sb
h0c/n_11895
h0c/n_12194
h0c/n_12614
h0c/n_6528
h0c/g64983_da
h0c/g64983_sb
h0c/n_4362
h0c/g64983_db
h0c/n_6234
h0c/g62655_da
h0c/g62655_db
h0c/g64973_da
h0c/g64973_sb
h0c/g64973_db
h0c/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__13__Q
h0c/g62655_sb
h0c/n_12112
h0c/n_12341
h0c/n_4432
h0c/g64853_db
h0c/g64853_da
h0c/g64853_sb
h0c/g63158_da
h0c/n_12009
h0c/g62963_db
h0c/n_4225
h0c/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__26__Q
h0c/n_5956
h0c/g65421_da
h0c/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__28__Q
h0c/g65421_sb
h0c/g62965_db
h0c/n_4226
h0c/g62965_sb
h0c/n_6526
h0c/g62525_da
h0c/g62525_db
h0c/wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__14__Q
h0c/g62525_sb
h0c/n_4371
h0c/g64972_da
h0c/g64972_db
h0c/g64972_sb
h0c/n_12868
h0c/g65043_sb
h0c/g65043_db
h0c/n_4326
h0c/g65334_sb
h0c/g62963_da
h0c/g62963_sb
h0c/n_5952
h0c/g62965_da
h0c/g64871_da
h0c/g64871_sb
h0c/n_12195
h0c/g65043_da
h0c/n_11993
h0c/g65335_sb
h0c/g64888_sb
h0c/n_11994
h0c/g65422_sb
h0c/g64993_sb
h0c/g65421_db
h0c/g64776_da
h0c/n_11984
h0c/n_16597
h0c/FE_OFN1171_n_4093
h0c/n_6490
h0c/g64871_db
h0c/g62539_db
h0c/n_4423
h0c/g65296_sb
h0c/n_3576
h0c/g65296_da
h0c/g65296_db
h0c/g65422_da
h0c/g65422_db
h0c/g64993_da
h0c/g64776_sb
h0c/n_12338
h0d/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__25__Q
h0d/n_10312
h0d/g57533_da
h0d/g57533_db
h0d/g57579_sb
h0d/g57579_db
h0d/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__26__Q
h0d/g58433_sb
h0d/n_11561
h0d/n_9006
h0d/g57533_sb
h0d/n_15589
h0d/g57579_da
h0d/n_9415
h0d/n_11173
h0d/g58433_da
h0d/n_10075
h0d/g57192_db
h0d/g58392_da
h0d/g58392_sb
h0d/g58396_db
h0d/g57538_sb
h0d/g58392_db
h0d/g58338_db
h0d/g58264_sb
h0d/g57549_da
h0d/n_9535
h0d/g57549_sb
h0d/n_11196
h0d/g57549_db
h0d/n_11260
h0d/g57477_da
h0d/g57477_db
h0d/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__7__Q
h0d/g58206_db
h0d/n_15595
h0d/n_9580
h0d/g58206_da
h0d/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_4__213
h0d/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__18__Q
h0d/n_11401
h0d/g57349_da
h0d/g57349_db
h0d/n_9005
h0d/g58396_da
h0d/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__2__Q
h0d/g58396_sb
h0d/g58264_db
h0d/g58264_da
h0d/n_9482
h0d/g57477_sb
h0d/n_15590
h0d/n_9303
h0d/g57349_sb
h0d/n_16842
h0d/g57538_db
h0d/g57538_da
h0d/g58338_da
h0d/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__7__Q
h0d/g58338_sb
h0d/g57466_sb
h0d/n_16836
h0d/n_15591
h0d/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__18__Q
h0d/g58115_da
h0d/g58115_sb
h0d/g58206_sb
h0d/g57043_db
h0d/n_10311
h0d/g58418_db
h0d/g58418_sb
h0d/g57923_db
h0d/n_11691
h0d/g57043_da
h0d/n_9887
h0d/g57923_da
h0d/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__2__Q
h0d/n_8998
h0d/g58418_da
h0d/n_15593
h0d/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__18__Q
h0d/n_11502
h0d/g57253_db
h0d/g57253_da
h0d/n_9678
h0d/g57253_sb
h0d/g57051_da
h0d/n_9132
h0d/g57051_sb
h0d/n_10509
h0d/g57051_db
h0d/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__25__Q
h0d/g57923_sb
h0d/n_11684
h0d/g57043_sb
h0d/n_10081
h0d/g57466_db
h0d/g57212_db
h0d/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__12__Q
h0d/n_10343
h0d/g57917_sb
h0d/g57466_da
h0d/g57037_sb
h0d/n_15586
h0d/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__12__Q
h0d/n_10515
h0d/g58115_db
h0d/n_16843
h0d/n_10439
h0d/g57212_da
h0d/g58072_db
h0d/n_9135
h0d/g57917_da
h0d/g57917_db
h0d/g58451_da
h0d/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__12__Q
h0d/g58451_sb
h0d/g57037_da
h0d/g57037_db
h0d/g57564_sb
h0d/g57564_db
h0d/n_15560
h0d/g58085_sb
h0d/g57931_da
h0d/g57931_db
h0d/g57931_sb
h0d/n_9084
h0d/g58085_da
h0d/g58085_db
h0d/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__25__Q
h0d/g57226_sb
h0d/n_10434
h0d/n_9087
h0d/g57212_sb
h0d/g58451_db
h0d/g57226_da
h0d/g57226_db
h0d/n_9328
h0d/n_9325
h0d/g58072_da
h0d/n_9280
h0d/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__25__Q
h0d/FE_OCPN1935_n_15566
h0d/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__25__Q
h0d/n_8991
h0d/g58432_sb
h0d/n_10297
h0d/g57578_da
h0d/n_8995
h0d/g57578_sb
h0d/g57066_da
h0d/n_9870
h0d/g57066_sb
h0d/g57943_sb
h0d/g57943_da
h0d/g57218_da
h0d/n_9716
h0d/g57218_sb
h0d/g58078_da
h0d/g58078_sb
h0d/n_10084
h0d/n_9283
h0d/g58072_sb
h0d/n_10451
h0d/g57177_da
h0d/g57177_db
h0d/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__12__Q
h0d/FE_OCP_RBN2066_n_16572
h0d/g57564_da
h0d/g58432_da
h0d/g58432_db
h0d/n_11724
h0d/g57943_db
h0d/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__7__Q
h0d/g58078_db
h0d/g58058_da
h0d/n_9095
h0d/g58042_da
h0d/g58042_db
h0d/g57191_db
h0d/g58054_db
h0d/n_10447
h0d/g57191_da
h0d/n_10292
h0d/g57578_db
h0d/FE_OFN578_n_9904
h0d/g58444_da
h0d/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__7__Q
h0d/g58444_sb
h0d/n_11676
h0d/g57066_db
h0d/n_10547
h0d/n_11538
h0d/n_15584
h0d/g57196_da
h0d/g58058_db
h0d/g57196_sb
h0d/g57177_sb
h0d/FE_OCP_RBN2068_n_16572
h0d/n_16837
h0d/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__7__Q
h0d/n_9409
h0d/g58444_db
h0d/g57241_db
h0d/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__12__Q
h0d/g57344_db
h0d/g58201_db
h0d/n_9091
h0d/n_12130
h0d/n_11718
h0d/g58201_da
h0d/g58201_sb
h0d/g58054_da
h0d/FE_OCPN1878_n_9991
h0d/n_9092
h0d/g57191_sb
h0d/g58214_da
h0d/g58214_sb
h0d/FE_OCP_RBN2067_n_16572
h0d/n_15585
h0d/n_15562
h0d/n_9962
h0d/n_11161
h0d/g57593_da
h0d/g57593_db
h0d/g57593_sb
h0d/n_9305
h0d/g58097_da
h0d/g58097_sb
h0d/g58097_db
h0d/g58135_da
h0d/n_10391
h0d/g57344_da
h0d/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__25__Q
h0d/n_9055
h0d/g57344_sb
h0d/n_10386
h0d/g58214_db
h0d/g57357_db
h0d/g57357_da
h0d/n_9052
h0d/g57357_sb
h0d/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__7__Q
h0d/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__7__Q
h0d/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_6__252
h0d/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_7__291
h0d/g57206_db
h0d/n_11551
h0d/n_10889
h0d/g57206_da
h0d/g58065_db
h0d/g57206_sb
h0d/g58065_da
h0d/g58065_sb
h0d/n_9727
h0d/n_11229
h0d/g58135_db
h0d/n_9661
h0d/g57273_sb
h0d/n_10864
h0d/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__7__Q
h0d/g57273_da
h0d/g57273_db
h0d/n_11482
h0d/g58007_da
h0d/g58007_sb
h0d/g58226_db
h0d/g58226_da
h0d/g58226_sb
h0d/g57369_sb
h0d/n_9563
h0d/g57369_da
h0d/n_11381
h0d/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__18__Q
h0d/n_11571
h0d/g57183_sb
h0d/n_15569
h0d/g57183_db
h0d/g57183_da
h0d/n_9742
h0d/g58047_db
h0d/g58047_da
h0d/g58047_sb
h0d/g58426_sb
h0d/g57077_db
h0d/g58007_db
h0d/n_11645
h0d/n_9787
h0d/g57101_da
h0d/g57101_sb
h0d/g57101_db
h0d/g58368_db
h0d/n_9458
h0d/g58368_da
h0d/g58368_sb
h0d/g57509_sb
h0d/g57369_db
h0d/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__3__Q
h0d/g57509_da
h0d/g57509_db
h0d/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__3__Q
h0d/n_11647
h0d/g57971_db
h0d/n_9829
h0d/g57971_da
h0d/g57100_da
h0d/g57100_sb
h0d/g57100_db
h0d/g57971_sb
h0d/g58147_da
h0d/g58147_sb
h0d/n_10193
h0d/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__13__Q
h0d/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__13__Q
h0d/g58422_sb
h0d/g58422_da
h0d/n_11187
h0d/g57565_da
h0d/g57565_db
h0d/g58422_db
h0d/n_9425
h0d/g58017_da
h0d/g58017_sb
h0d/g57565_sb
h0d/n_11230
h0d/n_9775
h0d/g58017_db
h0d/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__18__Q
h0d/g57148_da
h0d/g57148_sb
h0d/n_11602
h0d/g57148_db
h0d/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__18__Q
h0d/n_11468
h0d/g57285_sb
h0d/g57285_db
h0d/g57285_da
h0d/g58147_db
h0d/n_9647
h0d/g57948_sb
h0d/g58043_db
h0d/n_11577
h0d/g57178_da
h0d/g57178_db
h0d/g58043_da
h0d/g58043_sb
h0d/n_9746
h0d/g57178_sb
h0d/g58022_da
h0d/g58022_sb
h0d/g58022_db
h0d/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__22__Q
h0d/n_10463
h0d/g57153_da
h0d/g57153_db
h0d/g57115_db
h0d/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__18__Q
h0d/n_11631
h0d/g57115_da
h0d/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__18__Q
h0d/n_11431
h0d/g57320_db
h0d/n_9466
h0d/g58356_da
h0d/g58356_db
h0d/g58355_db
h0d/n_9101
h0d/g57153_sb
h0d/g57985_db
h0d/g57320_da
h0d/g58356_sb
h0d/n_9109
h0d/g57991_da
h0d/g57991_db
h0d/g57117_sb
h0d/g57991_sb
h0d/g58026_da
h0d/g58026_sb
h0d/n_9813
h0d/g57115_sb
h0d/g57158_sb
h0d/g57158_db
h0d/g58177_sb
h0d/n_9612
h0d/g58177_da
h0d/g58177_db
h0d/g58023_sb
h0d/n_11241
h0d/g57496_da
h0d/g57496_db
h0d/g57496_sb
h0d/n_9763
h0d/g58026_db
h0d/g57985_sb
h0d/g57985_da
h0d/n_11592
h0d/g57158_da
h0d/g57320_sb
h0d/g58012_db
h0d/g58012_da
h0d/g58012_sb
h0d/g58023_da
h0d/n_9767
h0d/g57155_sb
h1d/g58408_da
h1d/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__9__Q
h1d/g58408_sb
h1d/n_9432
h1d/g58408_db
h1d/g57551_sb
h1d/g58383_db
h1d/g57551_db
h1d/g57551_da
h1d/g58314_db
h1d/g58340_db
h1d/g58340_da
h1d/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__9__Q
h1d/g58340_sb
h1d/n_11193
h1d/g57479_da
h1d/n_9480
h1d/g57479_sb
h1d/n_11258
h1d/g57479_db
h1d/n_9491
h1d/g58322_db
h1d/g58309_db
h1d/n_11715
h1d/g58309_sb
h1d/g58309_da
h1d/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__11__Q
h1d/g57461_sb
h1d/n_9501
h1d/g57446_da
h1d/g57446_sb
h1d/g57532_da
h1d/n_9441
h1d/g58391_da
h1d/g58391_sb
h1d/g58391_db
h1d/g58377_sb
h1d/n_9452
h1d/g58377_da
h1d/g58377_db
h1d/n_11286
h1d/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__11__Q
h1d/g57446_db
h1d/n_11209
h1d/n_10994
h1d/FE_RN_186_0
h1d/g57939_da
h1d/g57939_sb
h1d/g57518_da
h1d/g57518_sb
h1d/n_11222
h1d/g57518_db
h1d/g57062_db
h1d/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__3__Q
h1d/g57036_da
h1d/n_9893
h1d/g57036_sb
h1d/g57916_sb
h1d/n_9871
h1d/g57939_db
h1d/g57062_sb
h1d/n_11677
h1d/g57062_da
h1d/n_11696
h1d/g57036_db
h1d/g57916_db
h1d/g57916_da
h1d/g58093_sb
h1d/g58093_da
h1d/g58093_db
h1d/g57237_sb
h1d/g58108_sb
h1d/n_9704
h1d/n_9662
h1d/g57269_sb
h1d/g57246_sb
h1d/g58108_da
h1d/n_9685
h1d/g58108_db
h1d/g58131_da
h1d/g58131_sb
h1d/g58131_db
h1d/g57246_db
h1d/n_11510
h1d/FE_RN_187_0
h1d/g57945_db
h1d/g57945_sb
h1d/n_10855
h1d/g57945_da
h1d/g57068_db
h1d/g57068_da
h1d/n_9867
h1d/g57246_da
h1d/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__3__Q
h1d/g57365_db
h1d/g57342_da
h1d/g58222_db
h1d/n_9564
h1d/g58222_da
h1d/g58222_sb
h1d/g57365_da
h1d/g57365_sb
h1d/n_11382
h1d/g58098_db
h1d/n_9702
h1d/g58098_da
h1d/g57243_sb
h1d/n_9585
h1d/g58114_da
h1d/g58114_sb
h1d/g58114_db
h1d/n_9680
h1d/g57252_sb
h1d/g58098_sb
h1d/g57252_da
h1d/g57252_db
h1d/n_11503
h1d/g58122_da
h1d/g58122_sb
h1d/g58213_sb
h1d/g58122_db
h1d/n_9670
h1d/g58205_sb
h1d/g57260_da
h1d/g57260_sb
h1d/g57260_db
h1d/g57348_db
h1d/n_11493
h1d/g58171_da
h1d/g58171_sb
h1d/g58205_da
h1d/g58205_db
h1d/n_9582
h1d/g58197_sb
h1d/g57348_da
h1d/g57348_sb
h1d/n_11402
h1d/n_9655
h1d/g57278_sb
h1d/g58197_db
h1d/g58197_da
h1d/n_9589
h1d/g57339_db
h1d/g57339_sb
h1d/n_11413
h1d/g57339_da
h1d/g57307_sb
h1d/g58140_da
h1d/g58140_sb
h1d/g57979_sb
h1d/g58168_sb
h1d/g57979_da
h1d/g58168_da
h1d/n_9623
h1d/g58168_db
h1d/g57106_sb
h1d/g57307_db
h1d/n_11443
h1d/g57307_da
h1d/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__11__Q
h1d/n_11639
h1d/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__11__Q
h1d/g57979_db
h1d/n_9820
h1d/g57106_da
h1d/g57141_sb
h1d/n_11607
h1d/g57141_da
h1d/g57141_db
h1d/g57106_db
h1d/g58010_sb
h1d/g58010_db
h1d/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__9__Q
h1d/wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__9__Q
h1d/g58038_sb
h1d/n_9783
h1d/g58010_da
h1d/n_9751
h1d/g58038_da
h1d/g58038_db
h1d/g57173_sb
h1d/g57173_da
h1d/n_11583
h1d/g57173_db
h1d/g58006_db
h1d/g58006_da
h1d/g58006_sb
h1d/g57138_da
h1d/n_9788
h1d/g57138_sb
h1d/n_11611
h1d/g57138_db
h1d/g58154_da
h1d/g58154_sb
h6/n_13715
h6/n_13716
h6/g57790_sb
h6/g67052_da
h6/g67052_sb
h6/FE_RN_329_0
h6/parity_checker_pci_perr_en_reg
h6/parity_checker_perr_sampled
h6/FE_RN_330_0
h6/g57790_da
h6/n_2254
h6/g67070_db
h6/g63215_p
h6/n_2249
h6/g57790_db
h6/n_14386
h6/n_13332
h6/n_13333
h6/g67070_da
h6/g64385_p
h6/n_1439
h6/n_2963
h6/FE_RN_304_0
h6/FE_RN_280_0
h6/n_7093
h6/FE_RN_306_0
h6/FE_RN_279_0
h6/n_13918
h6/FE_RN_149_0
h6/g53726_p
h6/g67070_sb
h6/FE_RN_305_0
h6/n_4699
h6/n_13758
h6/n_14765
h6/FE_RN_147_0
h6/FE_RN_148_0
h6/n_13335
h6/g54038_da
h6/g66014_p
h6/n_673
h6/g67146_p
h6/FE_RN_146_0
h6/g59782_p
h6/parchk_pci_perr_out_in
h6/n_14662
h6/parity_checker_check_perr
h6/parity_checker_check_perr_reg_Q
h6/g54038_sb
h6/g65945_sb
h6/g65945_da
h6/n_2576
h6/g65945_db
h6/FE_RN_144_0
h6/FE_RN_145_0
h6/output_backup_perr_out_reg_Q
h6/pci_target_unit_del_sync_addr_in_215
h6/FE_OFN1835_n_2678
h6/FE_OFN744_n_2678
h6/n_14624
h6/out_bckp_perr_en_out
h6/configuration_pci_err_data_505
h6/configuration_pci_err_addr_474
h6/pci_target_unit_pci_target_if_norm_address_reg_8__Q
h6/n_2611
h6/pci_target_unit_del_sync_addr_in_211
h6/FE_OFN1836_n_2678
h6/g66397_sb
h6/g66959_p
h6/pci_target_unit_pcit_if_strd_addr_in_697
h6/n_14572
h6/g66397_db
h6/n_2546
h6/g66397_da
h6/g65227_da
h6/g65227_sb
h6/n_722
h6/n_658
h6/g66934_p
h6/n_5662
h6/g60659_db
h6/g60659_da
h6/g65227_db
h6/g65928_sb
h6/g65928_da
h6/n_2507
h6/n_2660
h6/n_623
h6/g66947_p
h6/n_2583
h6/g65928_db
h6/pci_target_unit_del_sync_addr_in_229
h6/n_2667
h6/g65220_db
h6/g65220_da
h6/g65220_sb
h6/g66406_sb
h6/g65925_sb
h6/g65925_da
h6/g65231_db
h6/g65231_sb
h6/g66421_sb
h6/g65218_db
h6/n_2669
h6/g65218_da
h6/g65218_sb
h6/n_2586
h6/g65925_db
h6/n_2656
h6/g65231_da
h6/g65864_sb
h6/n_5656
h6/n_5664
h6/g65229_sb
h6/g65229_da
h6/pci_target_unit_del_sync_addr_in_216
h6/g66953_p
h6/g65864_da
h6/g60663_da
h6/g60663_db
h6/g60632_db
h6/g60657_db
h6/g65229_db
h6/n_2658
h6/g65864_db
h6/n_2593
h6/g67057_da
h6/g67054_sb
h6/n_1685
h6/n_5704
h6/g66405_db
h6/g66405_sb
h6/g66405_da
h6/g67057_db
h6/g67054_da
h6/g60632_da
h6/g67094_da
h6/n_613
h6/n_624
h6/n_2534
h6/g66937_p
h6/n_5654
h6/g60665_db
h6/n_5707
h6/g67054_db
h6/g60666_sb
h6/g65948_sb
h6/g52638_sb
h6/g52638_da
h6/g60665_da
h6/g60630_db
h6/g52649_da
h6/g52649_sb
h6/g65948_da
h6/g65219_db
h6/g52652_sb
h6/g52649_db
h6/g65948_db
h6/n_2668
h6/g65219_da
h6/g52638_db
h6/g60665_sb
h6/g60663_sb
h6/g52646_sb
h6/g52639_sb
h6/g52626_sb
h6/g65219_sb
h6/n_14645
h6/g60632_sb
h7
--pins(158)
FE_OFN1038_g64577_p
use :  
dir : o
shape : 
(3650,53490):(3750,54000) : 1
FE_OFN1047_g64577_p
use : �
dir : o
shape : 
(15250,53490):(15350,54000) : 1
FE_OFN1052_g64577_p
use :  
dir : o
shape : 
(0,33975):(255,34175) : 2
FE_OFN1057_g64577_p
use :  
dir : o
shape : 
(17650,53490):(17750,54000) : 1
FE_OFN1058_g64577_p
use :  
dir : o
shape : 
(5450,53490):(5550,54000) : 1
g62724_db
use :  
dir : o
shape : 
(0,32625):(510,32725) : 2
g62724_sb
use :  
dir : o
shape : 
(0,34825):(510,34925) : 2
g62776_sb
use :  
dir : o
shape : 
(8050,53490):(8150,54000) : 1
g62799_db
use :  
dir : o
shape : 
(2050,53490):(2150,54000) : 1
g62805_da
use :  
dir : o
shape : 
(5650,53490):(5750,54000) : 1
g62806_da
use :  
dir : o
shape : 
(30450,53490):(30550,54000) : 1
g62813_db
use :  
dir : o
shape : 
(3050,53490):(3150,54000) : 1
g62817_da
use :  
dir : o
shape : 
(1850,53490):(1950,54000) : 1
g62826_db
use :  
dir : o
shape : 
(0,24225):(510,24325) : 2
g63015_da
use :  
dir : o
shape : 
(24450,53490):(24550,54000) : 1
g63072_sb
use :  
dir : o
shape : 
(8250,53490):(8350,54000) : 1
g63105_db
use :  
dir : o
shape : 
(3850,53490):(3950,54000) : 1
g64152_sb
use :  
dir : o
shape : 
(0,45025):(510,45125) : 2
g64158_da
use :  
dir : o
shape : 
(0,30625):(510,30725) : 2
g64184_da
use :  
dir : o
shape : 
(0,42025):(510,42125) : 2
g64211_db
use :  
dir : o
shape : 
(3250,53490):(3350,54000) : 1
g64235_da
use :  
dir : o
shape : 
(0,44025):(510,44125) : 2
g64235_db
use :  
dir : o
shape : 
(0,45225):(510,45325) : 2
g64273_da
use :  
dir : o
shape : 
(14850,53490):(14950,54000) : 1
g64273_db
use :  
dir : o
shape : 
(15450,53490):(15550,54000) : 1
g64313_da
use :  
dir : o
shape : 
(7050,53490):(7150,54000) : 1
g64313_db
use :  
dir : o
shape : 
(0,45425):(510,45525) : 2
n_14060
use :  
dir : o
shape : 
(0,42625):(510,42725) : 2
n_14091
use :  
dir : o
shape : 
(0,45625):(510,45725) : 2
n_14092
use :  
dir : o
shape : 
(3450,53490):(3550,54000) : 1
n_14216
use :  
dir : o
shape : 
(0,38225):(510,38325) : 2
n_14596
use :  
dir : o
shape : 
(0,45825):(510,45925) : 2
n_14603
use :  
dir : o
shape : 
(27450,53490):(27550,54000) : 1
n_14608
use :  
dir : o
shape : 
(22050,53490):(22150,54000) : 1
n_14610
use :  
dir : o
shape : 
(26250,53490):(26350,54000) : 1
n_14611
use :  
dir : o
shape : 
(0,32825):(510,32925) : 2
n_16247
use :  
dir : o
shape : 
(21850,53490):(21950,54000) : 1
n_16252
use :  
dir : o
shape : 
(21650,53490):(21750,54000) : 1
n_3825
use :  
dir : o
shape : 
(6450,53490):(6550,54000) : 1
n_3938
use :  
dir : o
shape : 
(19450,53490):(19550,54000) : 1
n_3977
use :  
dir : o
shape : 
(0,26425):(510,26525) : 2
n_3983
use :  
dir : o
shape : 
(0,46025):(510,46125) : 2
n_4010
use :  
dir : o
shape : 
(0,47025):(510,47125) : 2
n_4077
use :  
dir : o
shape : 
(0,35025):(510,35125) : 2
n_5012
use :  
dir : o
shape : 
(4650,53490):(4750,54000) : 1
n_5136
use :  
dir : o
shape : 
(23450,53490):(23550,54000) : 1
n_5376
use :  
dir : o
shape : 
(0,46225):(510,46325) : 2
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__28__Q
use :  
dir : o
shape : 
(15850,53490):(15950,54000) : 1
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__28__Q
use :  
dir : o
shape : 
(8450,53490):(8550,54000) : 1
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__15__Q
use :  
dir : o
shape : 
(5050,53490):(5150,54000) : 3
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__18__Q
use :  
dir : o
shape : 
(0,43825):(510,43925) : 2
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__15__Q
use :  
dir : o
shape : 
(0,40225):(510,40325) : 2
pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_51
use :  
dir : o
shape : 
(99050,53490):(99150,54000) : 1
pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_63
use :  
dir : o
shape : 
(73850,53490):(73950,54000) : 1
FE_OCP_RBN2037_FE_OCPN2000_n_13743
use :  
dir : i
shape : 
(15650,53490):(15750,54000) : 1
FE_OCP_RBN2086_FE_OFN1756_n_13997
use :  
dir : i
shape : 
(32600,53745):(32800,54000) : 3
FE_OFN1015_g64577_p
use :  
dir : i
shape : 
(11450,53490):(11550,54000) : 1
FE_OFN1027_g64577_p
use :  
dir : i
shape : 
(0,37775):(255,37975) : 2
FE_OFN1034_g64577_p
use :  
dir : i
shape : 
(11200,53745):(11400,54000) : 3
FE_OFN1043_g64577_p
use :  
dir : i
shape : 
(33650,53490):(33750,54000) : 1
FE_OFN1046_g64577_p
use :  
dir : i
shape : 
(34200,53745):(34400,54000) : 3
FE_OFN1054_g64577_p
use :  
dir : i
shape : 
(32200,53745):(32400,54000) : 3
FE_OFN1464_n_13736
use :  
dir : i
shape : 
(0,39775):(255,39975) : 2
FE_OFN1465_n_13736
use :  
dir : i
shape : 
(23050,53490):(23150,54000) : 1
FE_OFN1466_n_13736
use :  
dir : i
shape : 
(43400,53745):(43600,54000) : 3
FE_OFN1469_n_13741
use :  
dir : i
shape : 
(0,34625):(510,34725) : 2
FE_OFN1470_n_13741
use :  
dir : i
shape : 
(28250,53490):(28350,54000) : 1
FE_OFN1471_n_13741
use :  
dir : i
shape : 
(4050,53490):(4150,54000) : 1
FE_OFN1478_n_13995
use :  
dir : i
shape : 
(24050,53490):(24150,54000) : 1
FE_OFN1479_n_13995
use :  
dir : i
shape : 
(7850,53490):(7950,54000) : 1
FE_OFN1522_n_4730
use :  
dir : i
shape : 
(15800,53745):(16000,54000) : 3
FE_OFN1523_n_4730
use :  
dir : i
shape : 
(35400,53745):(35600,54000) : 3
FE_OFN1524_n_4730
use :  
dir : i
shape : 
(0,33175):(255,33375) : 2
FE_OFN1557_n_4732
use :  
dir : i
shape : 
(0,38575):(255,38775) : 2
FE_OFN1558_n_4732
use :  
dir : i
shape : 
(33400,53745):(33600,54000) : 3
FE_OFN1559_n_4732
use :  
dir : i
shape : 
(7650,53490):(7750,54000) : 1
FE_OFN1581_n_16657
use :  
dir : i
shape : 
(0,41575):(255,41775) : 2
FE_OFN1583_n_16657
use :  
dir : i
shape : 
(31800,53745):(32000,54000) : 3
FE_OFN1584_n_16657
use :  
dir : i
shape : 
(0,39375):(255,39575) : 2
FE_OFN1612_n_4740
use :  
dir : i
shape : 
(0,40575):(255,40775) : 2
FE_OFN1613_n_4740
use :  
dir : i
shape : 
(5250,53490):(5350,54000) : 1
FE_OFN1614_n_4740
use :  
dir : i
shape : 
(6250,53490):(6350,54000) : 1
FE_OFN1757_n_13997
use :  
dir : i
shape : 
(7250,53490):(7350,54000) : 1
FE_OFN1761_n_14054
use :  
dir : i
shape : 
(4250,53490):(4350,54000) : 1
FE_OFN1762_n_14054
use :  
dir : i
shape : 
(0,42975):(255,43175) : 2
FE_OFN1764_n_14054
use :  
dir : i
shape : 
(12050,53490):(12150,54000) : 1
FE_OFN1770_n_13800
use :  
dir : i
shape : 
(8850,53490):(8950,54000) : 1
FE_OFN1771_n_13800
use :  
dir : i
shape : 
(11650,53490):(11750,54000) : 1
FE_OFN1772_n_13800
use :  
dir : i
shape : 
(0,31625):(510,31725) : 2
FE_OFN1776_n_13971
use :  
dir : i
shape : 
(33800,53745):(34000,54000) : 3
FE_OFN1777_n_13971
use :  
dir : i
shape : 
(32450,53490):(32550,54000) : 1
FE_OFN854_n_4736
use :  
dir : i
shape : 
(15050,53490):(15150,54000) : 1
FE_OFN855_n_4736
use :  
dir : i
shape : 
(33000,53745):(33200,54000) : 3
FE_OFN859_n_4734
use :  
dir : i
shape : 
(6850,53490):(6950,54000) : 1
FE_OFN860_n_4734
use :  
dir : i
shape : 
(0,38975):(255,39175) : 2
FE_OFN868_n_4725
use :  
dir : i
shape : 
(0,28175):(255,28375) : 2
FE_OFN951_n_4725
use :  
dir : i
shape : 
(31050,53490):(31150,54000) : 1
FE_OFN952_n_4725
use :  
dir : i
shape : 
(0,37375):(255,37575) : 2
FE_OFN975_n_4727
use :  
dir : i
shape : 
(24200,53745):(24400,54000) : 3
FE_OFN976_n_4727
use :  
dir : i
shape : 
(43000,53745):(43200,54000) : 3
g62803_da
use :  
dir : i
shape : 
(2850,53490):(2950,54000) : 1
g62805_sb
use :  
dir : i
shape : 
(6050,53490):(6150,54000) : 1
g62862_sb
use :  
dir : i
shape : 
(4450,53490):(4550,54000) : 1
g63015_sb
use :  
dir : i
shape : 
(24850,53490):(24950,54000) : 1
g63057_sb
use :  
dir : i
shape : 
(22850,53490):(22950,54000) : 1
g63058_da
use :  
dir : i
shape : 
(16450,53490):(16550,54000) : 1
g63072_da
use :  
dir : i
shape : 
(0,44825):(510,44925) : 2
g63122_da
use :  
dir : i
shape : 
(4850,53490):(4950,54000) : 1
g64078_da
use :  
dir : i
shape : 
(0,34425):(510,34525) : 2
g64158_sb
use :  
dir : i
shape : 
(0,30425):(510,30525) : 2
g64217_db
use :  
dir : i
shape : 
(30050,53490):(30150,54000) : 1
g64217_sb
use :  
dir : i
shape : 
(29250,53490):(29350,54000) : 1
g64296_db
use :  
dir : i
shape : 
(0,26225):(510,26325) : 2
ispd_clk
use :  
dir : i
shape : 
(0,43375):(255,43575) : 2
n_13891
use :  
dir : i
shape : 
(0,44625):(510,44725) : 2
n_13901
use :  
dir : i
shape : 
(0,31175):(255,31375) : 2
n_13987
use :  
dir : i
shape : 
(26850,53490):(26950,54000) : 1
n_13993
use :  
dir : i
shape : 
(19050,53490):(19150,54000) : 1
n_14001
use :  
dir : i
shape : 
(13650,53490):(13750,54000) : 1
n_14458
use :  
dir : i
shape : 
(27250,53490):(27350,54000) : 1
n_14472
use :  
dir : i
shape : 
(11850,53490):(11950,54000) : 1
n_14594
use :  
dir : i
shape : 
(100050,53490):(100150,54000) : 1
n_14956
use :  
dir : i
shape : 
(0,32425):(510,32525) : 2
n_16244
use :  
dir : i
shape : 
(22650,53490):(22750,54000) : 1
n_16621
use :  
dir : i
shape : 
(27650,53490):(27750,54000) : 1
n_3923
use :  
dir : i
shape : 
(14650,53490):(14750,54000) : 1
n_3958
use :  
dir : i
shape : 
(2250,53490):(2350,54000) : 1
n_4013
use :  
dir : i
shape : 
(0,44425):(510,44525) : 2
n_5351
use :  
dir : i
shape : 
(0,41025):(510,41125) : 2
n_5371
use :  
dir : i
shape : 
(7450,53490):(7550,54000) : 1
n_5388
use :  
dir : i
shape : 
(0,42425):(510,42525) : 2
pci_target_unit_fifos_pciw_addr_data_in_128
use :  
dir : i
shape : 
(6650,53490):(6750,54000) : 1
pci_target_unit_fifos_pciw_addr_data_in_132
use :  
dir : i
shape : 
(0,30825):(510,30925) : 2
pci_target_unit_fifos_pciw_addr_data_in_133
use :  
dir : i
shape : 
(32850,53490):(32950,54000) : 1
pci_target_unit_fifos_pciw_addr_data_in_134
use :  
dir : i
shape : 
(12250,53490):(12350,54000) : 1
pci_target_unit_fifos_pciw_addr_data_in_135
use :  
dir : i
shape : 
(35250,53490):(35350,54000) : 1
pci_target_unit_fifos_pciw_addr_data_in_136
use :  
dir : i
shape : 
(16850,53490):(16950,54000) : 1
pci_target_unit_fifos_pciw_addr_data_in_138
use :  
dir : i
shape : 
(26650,53490):(26750,54000) : 1
pci_target_unit_fifos_pciw_addr_data_in_141
use :  
dir : i
shape : 
(32250,53490):(32350,54000) : 1
pci_target_unit_fifos_pciw_addr_data_in_142
use :  
dir : i
shape : 
(0,41225):(510,41325) : 2
pci_target_unit_fifos_pciw_addr_data_in_148
use :  
dir : i
shape : 
(14450,53490):(14550,54000) : 1
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__13__Q
use :  
dir : i
shape : 
(24250,53490):(24350,54000) : 1
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__16__Q
use :  
dir : i
shape : 
(21450,53490):(21550,54000) : 1
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__13__Q
use :  
dir : i
shape : 
(23250,53490):(23350,54000) : 1
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__22__Q
use :  
dir : i
shape : 
(5850,53490):(5950,54000) : 1
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__8__Q
use :  
dir : i
shape : 
(0,46825):(510,46925) : 2
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__8__Q
use :  
dir : i
shape : 
(0,46625):(510,46725) : 2
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__12__Q
use :  
dir : i
shape : 
(0,30225):(510,30325) : 2
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__17__Q
use :  
dir : i
shape : 
(2450,53490):(2550,54000) : 1
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__28__Q
use :  
dir : i
shape : 
(0,44225):(510,44325) : 2
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__14__Q
use :  
dir : i
shape : 
(5050,53490):(5150,54000) : 1
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__21__Q
use :  
dir : i
shape : 
(28450,53490):(28550,54000) : 1
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__28__Q
use :  
dir : i
shape : 
(0,46425):(510,46525) : 2
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__13__Q
use :  
dir : i
shape : 
(0,33625):(510,33725) : 2
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__22__Q
use :  
dir : i
shape : 
(2650,53490):(2750,54000) : 1
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__12__Q
use :  
dir : i
shape : 
(0,29225):(510,29325) : 2
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__13__Q
use :  
dir : i
shape : 
(0,32225):(510,32325) : 2
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__15__Q
use :  
dir : i
shape : 
(0,42225):(510,42325) : 2
h8
--pins(268)
FE_OCP_RBN2089_FE_OFN1433_n_12042
use : _
dir : o
shape : 
(0,26900):(510,27000) : 2
FE_OCP_RBN2094_FE_OCPN1856_n_12030
use :  
dir : o
shape : 
(20050,49490):(20150,50000) : 1
FE_OFN1124_n_6935
use :  
dir : o
shape : 
(19450,49490):(19550,50000) : 1
FE_OFN1204_n_4097
use :  
dir : o
shape : 
(54000,49745):(54200,50000) : 3
FE_OFN1205_n_4097
use :  
dir : o
shape : 
(24850,49490):(24950,50000) : 1
FE_OFN1206_n_4097
use :  
dir : o
shape : 
(35400,49745):(35600,50000) : 3
FE_OFN1207_n_4097
use :  
dir : o
shape : 
(0,36850):(255,37050) : 2
FE_OFN1238_n_6436
use :  
dir : o
shape : 
(23450,49490):(23550,50000) : 1
FE_OFN1450_n_10780
use : z
dir : o
shape : 
(14250,49490):(14350,50000) : 1
FE_OFN1723_n_16317
use : z
dir : o
shape : 
(0,25500):(510,25600) : 2
FE_OFN647_n_4460
use : z
dir : o
shape : 
(32050,49490):(32150,50000) : 1
FE_OFN652_n_4417
use : z
dir : o
shape : 
(29200,0):(29400,255) : 3
FE_OFN658_n_4438
use : z
dir : o
shape : 
(22250,49490):(22350,50000) : 1
FE_RN_199_0
use : z
dir : o
shape : 
(17250,0):(17350,510) : 1
FE_RN_216_0
use : z
dir : o
shape : 
(21650,49490):(21750,50000) : 1
g54587_p
use : z
dir : o
shape : 
(26050,49490):(26150,50000) : 1
g62336_da
use :  
dir : o
shape : 
(19250,49490):(19350,50000) : 1
g62386_db
use :  
dir : o
shape : 
(16650,49490):(16750,50000) : 1
g62426_db
use :  
dir : o
shape : 
(23250,49490):(23350,50000) : 1
g62540_db
use :  
dir : o
shape : 
(21850,49490):(21950,50000) : 1
g62582_da
use :  
dir : o
shape : 
(0,26100):(510,26200) : 2
g62675_da
use :  
dir : o
shape : 
(22450,49490):(22550,50000) : 1
g62685_da
use :  
dir : o
shape : 
(49050,49490):(49150,50000) : 1
g62980_da
use :  
dir : o
shape : 
(70450,49490):(70550,50000) : 1
g62980_db
use :  
dir : o
shape : 
(71250,49490):(71350,50000) : 1
g64765_db
use :  
dir : o
shape : 
(18650,49490):(18750,50000) : 1
g64908_sb
use :  
dir : o
shape : 
(27850,49490):(27950,50000) : 1
g64949_da
use :  
dir : o
shape : 
(0,28100):(510,28200) : 2
g64974_db
use :  
dir : o
shape : 
(14850,49490):(14950,50000) : 1
g64993_db
use :  
dir : o
shape : 
(0,21700):(510,21800) : 2
g65004_db
use :  
dir : o
shape : 
(0,31100):(510,31200) : 2
g65047_sb
use :  
dir : o
shape : 
(18850,49490):(18950,50000) : 1
g65328_db
use :  
dir : o
shape : 
(15250,49490):(15350,50000) : 1
g65394_sb
use :  
dir : o
shape : 
(72850,49490):(72950,50000) : 1
n_11898
use :  
dir : o
shape : 
(16850,49490):(16950,50000) : 1
n_11899
use :  
dir : o
shape : 
(15650,49490):(15750,50000) : 1
n_11988
use :  
dir : o
shape : 
(0,26300):(510,26400) : 2
n_12002
use :  
dir : o
shape : 
(0,28300):(510,28400) : 2
n_12011
use :  
dir : o
shape : 
(0,30900):(510,31000) : 2
n_12041
use :  
dir : o
shape : 
(60050,49490):(60150,50000) : 1
n_12049
use :  
dir : o
shape : 
(70850,49490):(70950,50000) : 1
n_12052
use :  
dir : o
shape : 
(27450,49490):(27550,50000) : 1
n_12089
use :  
dir : o
shape : 
(0,31500):(510,31600) : 2
n_12102
use :  
dir : o
shape : 
(48050,49490):(48150,50000) : 1
n_12118
use :  
dir : o
shape : 
(56250,49490):(56350,50000) : 1
n_12196
use :  
dir : o
shape : 
(24250,49490):(24350,50000) : 1
n_12351
use :  
dir : o
shape : 
(15850,49490):(15950,50000) : 1
n_12406
use :  
dir : o
shape : 
(0,29700):(510,29800) : 2
n_12427
use :  
dir : o
shape : 
(43850,49490):(43950,50000) : 1
n_12449
use :  
dir : o
shape : 
(0,30700):(510,30800) : 2
n_12459
use :  
dir : o
shape : 
(0,26500):(510,26600) : 2
n_12473
use :  
dir : o
shape : 
(14650,49490):(14750,50000) : 1
n_12483
use :  
dir : o
shape : 
(40050,49490):(40150,50000) : 1
n_12492
use :  
dir : o
shape : 
(0,28500):(510,28600) : 2
n_12746
use :  
dir : o
shape : 
(38050,49490):(38150,50000) : 1
n_12749
use :  
dir : o
shape : 
(65250,49490):(65350,50000) : 1
n_12817
use :  
dir : o
shape : 
(47850,49490):(47950,50000) : 1
n_12886
use :  
dir : o
shape : 
(0,30500):(510,30600) : 2
n_12934
use :  
dir : o
shape : 
(48250,49490):(48350,50000) : 1
n_13128
use :  
dir : o
shape : 
(0,26700):(510,26800) : 2
n_13139
use :  
dir : o
shape : 
(17050,49490):(17150,50000) : 1
n_14311
use :  
dir : o
shape : 
(28050,49490):(28150,50000) : 1
n_14314
use :  
dir : o
shape : 
(28650,49490):(28750,50000) : 1
n_14381
use :  
dir : o
shape : 
(25450,49490):(25550,50000) : 1
n_16409
use :  
dir : o
shape : 
(62250,49490):(62350,50000) : 1
n_3744
use :  
dir : o
shape : 
(38600,49745):(38800,50000) : 3
n_3749
use :  
dir : o
shape : 
(20850,49490):(20950,50000) : 1
n_3761
use :  
dir : o
shape : 
(23650,49490):(23750,50000) : 1
n_4473
use :  
dir : o
shape : 
(17250,49490):(17350,50000) : 1
n_4478
use :  
dir : o
shape : 
(32450,49490):(32550,50000) : 1
n_5975
use :  
dir : o
shape : 
(16050,49490):(16150,50000) : 1
n_6231
use :  
dir : o
shape : 
(27850,0):(27950,510) : 1
n_6348
use :  
dir : o
shape : 
(20450,49490):(20550,50000) : 3
n_6935
use :  
dir : o
shape : 
(23850,49490):(23950,50000) : 1
parchk_pci_ad_out_in_1179
use :  
dir : o
shape : 
(36250,49490):(36350,50000) : 1
parchk_pci_ad_out_in_1181
use :  
dir : o
shape : 
(25250,49490):(25350,50000) : 1
parchk_pci_ad_out_in_1182
use :  
dir : o
shape : 
(39050,49490):(39150,50000) : 1
wbs_wbb3_2_wbb2_dat_o_i_105
use :  
dir : o
shape : 
(14850,0):(14950,510) : 1
wbs_wbb3_2_wbb2_dat_o_i_116
use :  
dir : o
shape : 
(18850,0):(18950,510) : 1
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__18__Q
use :  
dir : o
shape : 
(22650,49490):(22750,50000) : 1
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__37__Q
use :  
dir : o
shape : 
(35050,49490):(35150,50000) : 1
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__11__Q
use :  
dir : o
shape : 
(62850,49490):(62950,50000) : 1
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__26__Q
use :  
dir : o
shape : 
(29250,49490):(29350,50000) : 1
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__12__Q
use :  
dir : o
shape : 
(19050,49490):(19150,50000) : 1
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__6__Q
use :  
dir : o
shape : 
(14450,49490):(14550,50000) : 1
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__25__Q
use :  
dir : o
shape : 
(20450,49490):(20550,50000) : 1
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__26__Q
use :  
dir : o
shape : 
(34850,49490):(34950,50000) : 1
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__28__Q
use :  
dir : o
shape : 
(0,31700):(510,31800) : 2
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__28__Q
use :  
dir : o
shape : 
(0,19900):(510,20000) : 2
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__24__Q
use :  
dir : o
shape : 
(30650,49490):(30750,50000) : 1
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__5__Q
use :  
dir : o
shape : 
(45450,49490):(45550,50000) : 1
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__8__Q
use :  
dir : o
shape : 
(0,23500):(510,23600) : 2
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__11__Q
use :  
dir : o
shape : 
(40250,49490):(40350,50000) : 1
FE_OCPN1856_n_12030
use :  
dir : i
shape : 
(20650,49490):(20750,50000) : 1
FE_OCPN1857_n_12030
use :  
dir : i
shape : 
(0,29300):(510,29400) : 2
FE_OCPN1885_FE_OFN1454_n_12028
use :  
dir : i
shape : 
(64400,49745):(64600,50000) : 3
FE_OFN1120_n_6935
use :  
dir : i
shape : 
(69600,49745):(69800,50000) : 3
FE_OFN1127_n_4090
use :  
dir : i
shape : 
(24050,49490):(24150,50000) : 1
FE_OFN1128_n_4090
use :  
dir : i
shape : 
(0,19450):(255,19650) : 2
FE_OFN1132_n_6356
use :  
dir : i
shape : 
(52800,49745):(53000,50000) : 3
FE_OFN1135_n_4151
use :  
dir : i
shape : 
(0,31450):(255,31650) : 4
FE_OFN1140_n_6886
use :  
dir : i
shape : 
(60850,49490):(60950,50000) : 1
FE_OFN1147_n_6391
use :  
dir : i
shape : 
(0,20250):(255,20450) : 2
FE_OFN1148_n_6391
use :  
dir : i
shape : 
(0,40450):(255,40650) : 2
FE_OFN1156_n_6391
use :  
dir : i
shape : 
(71800,49745):(72000,50000) : 3
FE_OFN1159_n_6391
use :  
dir : i
shape : 
(54800,0):(55000,255) : 3
FE_OFN1162_n_6391
use :  
dir : i
shape : 
(38200,49745):(38400,50000) : 3
FE_OFN1167_n_4092
use :  
dir : i
shape : 
(23200,0):(23400,255) : 3
FE_OFN1174_n_4093
use :  
dir : i
shape : 
(0,16650):(255,16850) : 2
FE_OFN1177_n_4143
use :  
dir : i
shape : 
(38650,49490):(38750,50000) : 1
FE_OFN1184_n_4143
use :  
dir : i
shape : 
(0,38850):(255,39050) : 2
FE_OFN1185_n_4143
use :  
dir : i
shape : 
(37800,49745):(38000,50000) : 3
FE_OFN1189_n_4095
use :  
dir : i
shape : 
(36000,0):(36200,255) : 3
FE_OFN1190_n_4095
use :  
dir : i
shape : 
(56600,49745):(56800,50000) : 3
FE_OFN1193_n_4095
use :  
dir : i
shape : 
(33400,0):(33600,255) : 3
FE_OFN1198_n_4096
use :  
dir : i
shape : 
(0,32850):(255,33050) : 2
FE_OFN119_n_12502
use :  
dir : i
shape : 
(0,31300):(510,31400) : 2
FE_OFN1213_n_4098
use :  
dir : i
shape : 
(40200,0):(40400,255) : 3
FE_OFN1225_n_6624
use :  
dir : i
shape : 
(0,38450):(255,38650) : 2
FE_OFN1226_n_6624
use :  
dir : i
shape : 
(39400,0):(39600,255) : 3
FE_OFN1231_n_6624
use :  
dir : i
shape : 
(36400,0):(36600,255) : 3
FE_OFN1233_n_6624
use :  
dir : i
shape : 
(59000,49745):(59200,50000) : 3
FE_OFN1235_n_6436
use :  
dir : i
shape : 
(25850,49490):(25950,50000) : 1
FE_OFN130_n_12104
use :  
dir : i
shape : 
(47450,49490):(47550,50000) : 1
FE_OFN1431_n_12104
use :  
dir : i
shape : 
(16250,49490):(16350,50000) : 1
FE_OFN1435_n_12042
use :  
dir : i
shape : 
(73000,49745):(73200,50000) : 3
FE_OFN1441_n_12502
use :  
dir : i
shape : 
(28450,49490):(28550,50000) : 1
FE_OFN1445_n_12502
use :  
dir : i
shape : 
(70800,49745):(71000,50000) : 3
FE_OFN1449_n_10780
use :  
dir : i
shape : 
(21250,49490):(21350,50000) : 1
FE_OFN1455_n_12028
use :  
dir : i
shape : 
(0,37250):(255,37450) : 2
FE_OFN1458_n_12306
use :  
dir : i
shape : 
(24450,49490):(24550,50000) : 1
FE_OFN1461_n_12306
use :  
dir : i
shape : 
(17850,49490):(17950,50000) : 1
FE_OFN1474_n_14995
use :  
dir : i
shape : 
(39250,49490):(39350,50000) : 1
FE_OFN1475_n_14995
use :  
dir : i
shape : 
(15050,49490):(15150,50000) : 1
FE_OFN1507_n_4460
use :  
dir : i
shape : 
(31450,49490):(31550,50000) : 1
FE_OFN1511_n_4460
use :  
dir : i
shape : 
(0,30050):(255,30250) : 2
FE_OFN1515_n_4677
use :  
dir : i
shape : 
(16200,0):(16400,255) : 3
FE_OFN1547_n_4501
use :  
dir : i
shape : 
(0,37650):(255,37850) : 2
FE_OFN1548_n_4501
use :  
dir : i
shape : 
(35250,49490):(35350,50000) : 1
FE_OFN1549_n_4501
use :  
dir : i
shape : 
(54600,49745):(54800,50000) : 3
FE_OFN1653_n_4868
use :  
dir : i
shape : 
(37400,49745):(37600,50000) : 3
FE_OFN1654_n_4868
use :  
dir : i
shape : 
(12600,49745):(12800,50000) : 3
FE_OFN1718_n_16317
use :  
dir : i
shape : 
(26450,49490):(26550,50000) : 1
FE_OFN1726_n_14987
use :  
dir : i
shape : 
(44050,49490):(44150,50000) : 1
FE_OFN1733_n_11019
use :  
dir : i
shape : 
(26250,0):(26350,510) : 1
FE_OFN1745_n_12086
use :  
dir : i
shape : 
(0,32500):(510,32600) : 2
FE_OFN1751_n_11027
use :  
dir : i
shape : 
(0,29500):(510,29600) : 4
FE_OFN1755_n_12681
use :  
dir : i
shape : 
(16650,0):(16750,510) : 1
FE_OFN1794_n_4508
use :  
dir : i
shape : 
(0,31050):(255,31250) : 4
FE_OFN1797_n_4508
use :  
dir : i
shape : 
(0,39850):(255,40050) : 2
FE_OFN1804_n_3741
use :  
dir : i
shape : 
(0,27450):(255,27650) : 2
FE_OFN1826_n_4490
use :  
dir : i
shape : 
(57000,49745):(57200,50000) : 3
FE_OFN325_g66125_p
use :  
dir : i
shape : 
(23050,49490):(23150,50000) : 1
FE_OFN589_n_4490
use :  
dir : i
shape : 
(53600,49745):(53800,50000) : 3
FE_OFN590_n_4490
use :  
dir : i
shape : 
(0,41050):(255,41250) : 2
FE_OFN591_n_4490
use :  
dir : i
shape : 
(39000,49745):(39200,50000) : 3
FE_OFN595_n_4409
use :  
dir : i
shape : 
(29200,49745):(29400,50000) : 3
FE_OFN596_n_4409
use :  
dir : i
shape : 
(0,28050):(255,28250) : 4
FE_OFN597_n_4409
use :  
dir : i
shape : 
(57400,49745):(57600,50000) : 3
FE_OFN599_n_4454
use :  
dir : i
shape : 
(36200,49745):(36400,50000) : 3
FE_OFN600_n_4454
use :  
dir : i
shape : 
(0,34450):(255,34650) : 2
FE_OFN607_n_4669
use :  
dir : i
shape : 
(35800,49745):(36000,50000) : 3
FE_OFN612_n_4497
use :  
dir : i
shape : 
(0,35450):(255,35650) : 2
FE_OFN613_n_4497
use :  
dir : i
shape : 
(69200,49745):(69400,50000) : 3
FE_OFN614_n_4497
use :  
dir : i
shape : 
(0,22050):(255,22250) : 2
FE_OFN626_n_4392
use :  
dir : i
shape : 
(20200,0):(20400,255) : 3
FE_OFN629_n_4495
use :  
dir : i
shape : 
(0,38050):(255,38250) : 2
FE_OFN631_n_4495
use :  
dir : i
shape : 
(0,23050):(255,23250) : 2
FE_OFN634_n_4505
use :  
dir : i
shape : 
(0,39450):(255,39650) : 2
FE_OFN635_n_4505
use :  
dir : i
shape : 
(72200,49745):(72400,50000) : 3
FE_OFN636_n_4505
use :  
dir : i
shape : 
(34200,49745):(34400,50000) : 3
FE_OFN649_n_4417
use :  
dir : i
shape : 
(27650,49490):(27750,50000) : 1
FE_OFN654_n_4438
use :  
dir : i
shape : 
(26250,49490):(26350,50000) : 1
FE_OFN656_n_4438
use :  
dir : i
shape : 
(35600,0):(35800,255) : 3
FE_OFN967_n_4655
use :  
dir : i
shape : 
(55000,49745):(55200,50000) : 3
FE_OFN968_n_4655
use :  
dir : i
shape : 
(35000,0):(35200,255) : 3
FE_RN_203_0
use :  
dir : i
shape : 
(17650,49490):(17750,50000) : 1
g62336_sb
use :  
dir : i
shape : 
(19850,49490):(19950,50000) : 1
g62345_da
use :  
dir : i
shape : 
(0,42500):(510,42600) : 2
g62362_db
use :  
dir : i
shape : 
(0,42300):(510,42400) : 2
g62362_sb
use :  
dir : i
shape : 
(21450,49490):(21550,50000) : 1
g62389_db
use :  
dir : i
shape : 
(33250,49490):(33350,50000) : 1
g62389_sb
use :  
dir : i
shape : 
(32250,49490):(32350,50000) : 1
g62410_db
use :  
dir : i
shape : 
(0,29500):(510,29600) : 2
g62485_sb
use :  
dir : i
shape : 
(24650,49490):(24750,50000) : 1
g62547_db
use :  
dir : i
shape : 
(47650,49490):(47750,50000) : 1
g62601_sb
use :  
dir : i
shape : 
(0,42100):(510,42200) : 2
g62911_db
use :  
dir : i
shape : 
(11050,49490):(11150,50000) : 3
g62923_db
use :  
dir : i
shape : 
(16450,49490):(16550,50000) : 1
g62923_sb
use :  
dir : i
shape : 
(11050,49490):(11150,50000) : 1
g62953_db
use :  
dir : i
shape : 
(10850,49490):(10950,50000) : 3
g62980_sb
use :  
dir : i
shape : 
(71050,49490):(71150,50000) : 1
g63183_da
use :  
dir : i
shape : 
(0,35900):(510,36000) : 2
g64800_sb
use :  
dir : i
shape : 
(42650,49490):(42750,50000) : 1
g64906_sb
use :  
dir : i
shape : 
(50850,49490):(50950,50000) : 1
g64907_sb
use :  
dir : i
shape : 
(56450,49490):(56550,50000) : 1
g64908_da
use :  
dir : i
shape : 
(25050,49490):(25150,50000) : 1
g64949_sb
use :  
dir : i
shape : 
(0,27900):(510,28000) : 2
g65335_da
use :  
dir : i
shape : 
(10850,49490):(10950,50000) : 1
g65351_sb
use :  
dir : i
shape : 
(73650,49490):(73750,50000) : 1
g65381_db
use :  
dir : i
shape : 
(29650,49490):(29750,50000) : 1
g65394_da
use :  
dir : i
shape : 
(72250,49490):(72350,50000) : 1
g65394_db
use :  
dir : i
shape : 
(72450,49490):(72550,50000) : 1
g66098_p
use :  
dir : i
shape : 
(31050,49490):(31150,50000) : 1
g66128_p
use :  
dir : i
shape : 
(21050,49490):(21150,50000) : 1
g66134_p
use :  
dir : i
shape : 
(10650,49490):(10750,50000) : 3
ispd_clk
use :  
dir : i
shape : 
(20250,49490):(20350,50000) : 1
n_12001
use :  
dir : i
shape : 
(0,26500):(510,26600) : 4
n_12010
use :  
dir : i
shape : 
(0,30650):(255,30850) : 4
n_12042
use :  
dir : i
shape : 
(10650,49490):(10750,50000) : 1
n_12105
use :  
dir : i
shape : 
(38450,49490):(38550,50000) : 1
n_12356
use :  
dir : i
shape : 
(0,33300):(510,33400) : 2
n_12403
use :  
dir : i
shape : 
(19250,0):(19350,510) : 1
n_12433
use :  
dir : i
shape : 
(49850,49490):(49950,50000) : 1
n_12458
use :  
dir : i
shape : 
(0,28500):(510,28600) : 4
n_12612
use :  
dir : i
shape : 
(0,25900):(510,26000) : 2
n_12645
use :  
dir : i
shape : 
(0,32100):(510,32200) : 4
n_12685
use :  
dir : i
shape : 
(62450,49490):(62550,50000) : 1
n_12695
use :  
dir : i
shape : 
(18450,49490):(18550,50000) : 1
n_12865
use :  
dir : i
shape : 
(0,32300):(510,32400) : 4
n_12866
use :  
dir : i
shape : 
(0,25700):(510,25800) : 2
n_13058
use :  
dir : i
shape : 
(10450,49490):(10550,50000) : 3
n_13144
use :  
dir : i
shape : 
(19850,0):(19950,510) : 1
n_13402
use :  
dir : i
shape : 
(16050,0):(16150,510) : 1
n_13760
use :  
dir : i
shape : 
(28250,49490):(28350,50000) : 1
n_14309
use :  
dir : i
shape : 
(40850,49490):(40950,50000) : 1
n_14313
use :  
dir : i
shape : 
(29050,49490):(29150,50000) : 1
n_14317
use :  
dir : i
shape : 
(36850,49490):(36950,50000) : 1
n_14353
use :  
dir : i
shape : 
(0,41900):(510,42000) : 2
n_156
use :  
dir : i
shape : 
(11250,49490):(11350,50000) : 1
n_3464
use :  
dir : i
shape : 
(12200,49745):(12400,50000) : 3
n_3752
use :  
dir : i
shape : 
(51000,49745):(51200,50000) : 3
n_3755
use :  
dir : i
shape : 
(56200,49745):(56400,50000) : 3
n_3770
use :  
dir : i
shape : 
(70000,49745):(70200,50000) : 3
n_3774
use :  
dir : i
shape : 
(72600,49745):(72800,50000) : 3
n_3777
use :  
dir : i
shape : 
(11800,49745):(12000,50000) : 3
n_3785
use :  
dir : i
shape : 
(18250,49490):(18350,50000) : 1
n_3792
use :  
dir : i
shape : 
(55400,49745):(55600,50000) : 3
n_4308
use :  
dir : i
shape : 
(0,31900):(510,32000) : 4
n_4357
use :  
dir : i
shape : 
(15050,0):(15150,510) : 1
n_4373
use :  
dir : i
shape : 
(17450,49490):(17550,50000) : 1
n_4442
use :  
dir : i
shape : 
(0,22450):(255,22650) : 2
n_4444
use :  
dir : i
shape : 
(49200,49745):(49400,50000) : 3
n_4450
use :  
dir : i
shape : 
(37000,49745):(37200,50000) : 3
n_4452
use :  
dir : i
shape : 
(36600,49745):(36800,50000) : 3
n_4465
use :  
dir : i
shape : 
(34200,0):(34400,255) : 3
n_4476
use :  
dir : i
shape : 
(34600,0):(34800,255) : 3
n_4479
use :  
dir : i
shape : 
(11400,49745):(11600,50000) : 3
n_4488
use :  
dir : i
shape : 
(55800,49745):(56000,50000) : 3
n_4493
use :  
dir : i
shape : 
(18000,0):(18200,255) : 3
n_4645
use :  
dir : i
shape : 
(0,32050):(255,32250) : 2
n_6189
use :  
dir : i
shape : 
(19650,49490):(19750,50000) : 1
n_6232
use :  
dir : i
shape : 
(53200,49745):(53400,50000) : 3
n_6287
use :  
dir : i
shape : 
(0,41450):(255,41650) : 2
n_6319
use :  
dir : i
shape : 
(30400,49745):(30600,50000) : 3
n_6388
use :  
dir : i
shape : 
(15850,0):(15950,510) : 1
n_6645
use :  
dir : i
shape : 
(13000,49745):(13200,50000) : 3
n_7631
use :  
dir : i
shape : 
(28850,49490):(28950,50000) : 1
n_7671
use :  
dir : i
shape : 
(25650,49490):(25750,50000) : 1
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__0__Q
use :  
dir : i
shape : 
(18050,49490):(18150,50000) : 1
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__29__Q
use :  
dir : i
shape : 
(22050,49490):(22150,50000) : 1
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__8__Q
use :  
dir : i
shape : 
(10450,49490):(10550,50000) : 1
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__12__Q
use :  
dir : i
shape : 
(15650,49490):(15750,50000) : 3
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__21__Q
use :  
dir : i
shape : 
(48850,49490):(48950,50000) : 1
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__29__Q
use :  
dir : i
shape : 
(22850,49490):(22950,50000) : 1
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__30__Q
use :  
dir : i
shape : 
(63450,49490):(63550,50000) : 1
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__16__Q
use :  
dir : i
shape : 
(70650,49490):(70750,50000) : 1
wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__14__Q
use :  
dir : i
shape : 
(0,21500):(510,21600) : 2
hh4
--pins(140)
FE_OCP_RBN2106_n_9155
use : ;
dir : o
shape : 
(352090,63750):(352600,63850) : 2
FE_OFN1262_n_8567
use :  
dir : o
shape : 
(352090,63950):(352600,64050) : 2
FE_OFN1316_n_8567
use :  
dir : o
shape : 
(182200,159745):(182400,160000) : 3
FE_OFN1334_n_9372
use :  
dir : o
shape : 
(352090,66150):(352600,66250) : 2
FE_OFN1336_n_9372
use :  
dir : o
shape : 
(352345,38900):(352600,39100) : 2
FE_OFN1337_n_9372
use : 9
dir : o
shape : 
(352345,39300):(352600,39500) : 2
FE_OFN1340_n_9372
use : �
dir : o
shape : 
(352345,64300):(352600,64500) : 2
FE_OFN1498_n_9864
use :  
dir : o
shape : 
(286450,0):(286550,510) : 1
FE_OFN1499_n_9864
use : �
dir : o
shape : 
(352345,64700):(352600,64900) : 2
FE_OFN1537_n_9428
use : Q
dir : o
shape : 
(171600,159745):(171800,160000) : 3
FE_OFN222_n_9844
use : \
dir : o
shape : 
(352345,13300):(352600,13500) : 2
FE_OFN248_n_9114
use : C
dir : o
shape : 
(352345,138700):(352600,138900) : 2
FE_OFN257_n_8969
use : 
dir : o
shape : 
(261850,159490):(261950,160000) : 1
FE_OFN448_n_10853
use : ?
dir : o
shape : 
(352090,65150):(352600,65250) : 2
FE_OFN523_n_9690
use : m
dir : o
shape : 
(289200,0):(289400,255) : 3
FE_OFN534_n_9864
use : P
dir : o
shape : 
(131800,0):(132000,255) : 3
FE_OFN566_n_9692
use :  
dir : o
shape : 
(352345,65500):(352600,65700) : 2
g57223_da
use :  
dir : o
shape : 
(202050,0):(202150,510) : 1
g57530_db
use :  
dir : o
shape : 
(95850,159490):(95950,160000) : 1
g57535_sb
use :  
dir : o
shape : 
(82850,0):(82950,510) : 1
g57913_db
use :  
dir : o
shape : 
(59050,0):(59150,510) : 1
g58063_sb
use :  
dir : o
shape : 
(24450,0):(24550,510) : 1
g58199_da
use :  
dir : o
shape : 
(128650,0):(128750,510) : 1
g58376_db
use :  
dir : o
shape : 
(126850,159490):(126950,160000) : 1
g58389_da
use :  
dir : o
shape : 
(105850,159490):(105950,160000) : 1
g58428_sb
use :  
dir : o
shape : 
(159050,159490):(159150,160000) : 1
g58439_db
use :  
dir : o
shape : 
(161050,159490):(161150,160000) : 1
g58439_sb
use :  
dir : o
shape : 
(164450,159490):(164550,160000) : 1
g58481_db
use :  
dir : o
shape : 
(278850,159490):(278950,160000) : 1
g58832_da
use :  
dir : o
shape : 
(266250,159490):(266350,160000) : 1
n_10185
use :  
dir : o
shape : 
(231050,0):(231150,510) : 1
n_10627
use :  
dir : o
shape : 
(257450,0):(257550,510) : 1
n_10753
use :  
dir : o
shape : 
(0,138350):(510,138450) : 2
n_11005
use : A
dir : o
shape : 
(265450,0):(265550,510) : 1
n_11236
use :  
dir : o
shape : 
(166850,0):(166950,510) : 1
n_11410
use :  
dir : o
shape : 
(321450,0):(321550,510) : 1
n_12573
use :  
dir : o
shape : 
(176650,0):(176750,510) : 1
n_12578
use : �
dir : o
shape : 
(278450,0):(278550,510) : 1
n_2933
use : Z
dir : o
shape : 
(352090,113350):(352600,113450) : 2
n_8714
use : �
dir : o
shape : 
(78650,159490):(78750,160000) : 1
n_8884
use :  
dir : o
shape : 
(223800,159745):(224000,160000) : 3
n_9228
use : �
dir : o
shape : 
(232250,159490):(232350,160000) : 1
n_9419
use : r
dir : o
shape : 
(98250,159490):(98350,160000) : 1
n_9440
use :  
dir : o
shape : 
(118250,0):(118350,510) : 1
wbu_sel_in_312
use : �
dir : o
shape : 
(238250,0):(238350,510) : 1
wishbone_slave_unit_del_sync_addr_out_reg_5__Q
use : �
dir : o
shape : 
(112850,159490):(112950,160000) : 1
wishbone_slave_unit_fifos_wbr_be_in_264
use :  
dir : o
shape : 
(352090,112950):(352600,113050) : 2
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__16__Q
use : �
dir : o
shape : 
(298450,0):(298550,510) : 1
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__31__Q
use :  
dir : o
shape : 
(352090,90150):(352600,90250) : 2
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__33__Q
use : 
dir : o
shape : 
(80450,159490):(80550,160000) : 1
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__10__Q
use :  
dir : o
shape : 
(275450,0):(275550,510) : 1
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__22__Q
use : N
dir : o
shape : 
(186450,0):(186550,510) : 1
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__20__Q
use :  
dir : o
shape : 
(0,89550):(510,89650) : 2
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__5__Q
use :  
dir : o
shape : 
(0,89350):(510,89450) : 2
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__27__Q
use :  
dir : o
shape : 
(220850,0):(220950,510) : 1
wishbone_slave_unit_pcim_if_wbw_addr_data_in_388
use : 
dir : o
shape : 
(352090,90350):(352600,90450) : 2
FE_OCPN1879_n_9991
use : �
dir : i
shape : 
(0,138550):(510,138650) : 2
FE_OCPN1936_n_15566
use : l
dir : i
shape : 
(257600,0):(257800,255) : 3
FE_OCP_RBN2104_n_9155
use : f
dir : i
shape : 
(352090,63550):(352600,63650) : 2
FE_OFN1251_n_16439
use : �
dir : i
shape : 
(267850,159490):(267950,160000) : 1
FE_OFN1253_n_8567
use : �
dir : i
shape : 
(352090,63350):(352600,63450) : 2
FE_OFN1282_n_8567
use : �
dir : i
shape : 
(179050,159490):(179150,160000) : 1
FE_OFN1285_n_8567
use : D
dir : i
shape : 
(0,112900):(255,113100) : 2
FE_OFN1287_n_8567
use : M
dir : i
shape : 
(211800,0):(212000,255) : 3
FE_OFN1289_n_8567
use :  
dir : i
shape : 
(331000,0):(331200,255) : 3
FE_OFN1296_n_8567
use :  
dir : i
shape : 
(88600,0):(88800,255) : 3
FE_OFN1298_n_8567
use :  
dir : i
shape : 
(65600,159745):(65800,160000) : 3
FE_OFN1308_n_8567
use :  
dir : i
shape : 
(95400,159745):(95600,160000) : 3
FE_OFN1315_n_8567
use :  
dir : i
shape : 
(133200,0):(133400,255) : 3
FE_OFN1341_n_9372
use :  
dir : i
shape : 
(269400,159745):(269600,160000) : 3
FE_OFN1377_n_10853
use :  
dir : i
shape : 
(352090,62950):(352600,63050) : 4
FE_OFN13_n_11877
use :  
dir : i
shape : 
(255200,0):(255400,255) : 3
FE_OFN1400_n_10566
use :  
dir : i
shape : 
(196450,0):(196550,510) : 1
FE_OFN1496_n_9864
use :  
dir : i
shape : 
(132050,0):(132150,510) : 1
FE_OFN1497_n_9864
use :  
dir : i
shape : 
(352090,62950):(352600,63050) : 2
FE_OFN1534_n_9428
use :  
dir : i
shape : 
(174050,159490):(174150,160000) : 1
FE_OFN1541_n_9502
use :  
dir : i
shape : 
(137850,159490):(137950,160000) : 1
FE_OFN1572_n_9477
use :  
dir : i
shape : 
(116200,159745):(116400,160000) : 3
FE_OFN1632_n_9862
use :  
dir : i
shape : 
(128000,159745):(128200,160000) : 3
FE_OFN1687_n_15534
use :  
dir : i
shape : 
(285850,0):(285950,510) : 1
FE_OFN1692_n_16992
use :  
dir : i
shape : 
(286250,0):(286350,510) : 1
FE_OFN1713_n_9320
use :  
dir : i
shape : 
(195850,0):(195950,510) : 1
FE_OFN1807_n_9899
use :  
dir : i
shape : 
(0,113900):(255,114100) : 2
FE_OFN199_n_9228
use :  
dir : i
shape : 
(161250,159490):(161350,160000) : 1
FE_OFN214_n_9856
use :  
dir : i
shape : 
(117400,0):(117600,255) : 3
FE_OFN220_n_9846
use :  
dir : i
shape : 
(128400,159745):(128600,160000) : 3
FE_OFN224_n_9122
use :  
dir : i
shape : 
(137400,159745):(137600,160000) : 3
FE_OFN233_n_9876
use :  
dir : i
shape : 
(108600,0):(108800,255) : 3
FE_OFN236_n_9834
use :  
dir : i
shape : 
(171200,159745):(171400,160000) : 3
FE_OFN498_n_9697
use :  
dir : i
shape : 
(196200,159745):(196400,160000) : 3
FE_OFN519_n_9690
use :  
dir : i
shape : 
(289450,0):(289550,510) : 1
FE_OFN548_n_9502
use :  
dir : i
shape : 
(152600,159745):(152800,160000) : 3
FE_OFN555_n_9902
use :  
dir : i
shape : 
(162200,0):(162400,255) : 3
FE_OFN559_n_9531
use :  
dir : i
shape : 
(109000,0):(109200,255) : 3
FE_OFN561_n_9692
use :  
dir : i
shape : 
(352090,63150):(352600,63250) : 2
FE_OFN571_n_9694
use :  
dir : i
shape : 
(165200,159745):(165400,160000) : 3
FE_OFN581_n_9904
use :  
dir : i
shape : 
(0,88900):(255,89100) : 2
g57041_da
use :  
dir : i
shape : 
(306250,0):(306350,510) : 1
g57341_db
use :  
dir : i
shape : 
(321050,0):(321150,510) : 1
g58063_da
use :  
dir : i
shape : 
(0,38950):(510,39050) : 2
g58082_db
use :  
dir : i
shape : 
(171250,0):(171350,510) : 1
g58361_da
use :  
dir : i
shape : 
(142650,0):(142750,510) : 1
g58389_sb
use :  
dir : i
shape : 
(106250,159490):(106350,160000) : 1
g58393_da
use :  
dir : i
shape : 
(118450,0):(118550,510) : 1
g58428_da
use :  
dir : i
shape : 
(98450,159490):(98550,160000) : 1
g58829_db
use :  
dir : i
shape : 
(210850,159490):(210950,160000) : 1
g59091_da
use :  
dir : i
shape : 
(78850,159490):(78950,160000) : 1
g59091_db
use :  
dir : i
shape : 
(79050,159490):(79150,160000) : 1
g63585_da
use :  
dir : i
shape : 
(244450,0):(244550,510) : 1
ispd_clk
use :  
dir : i
shape : 
(251000,0):(251200,255) : 3
n_10051
use :  
dir : i
shape : 
(160650,0):(160750,510) : 1
n_10054
use :  
dir : i
shape : 
(166050,0):(166150,510) : 1
n_10057
use :  
dir : i
shape : 
(165050,0):(165150,510) : 1
n_10314
use :  
dir : i
shape : 
(111450,159490):(111550,160000) : 1
n_10693
use :  
dir : i
shape : 
(0,138750):(510,138850) : 2
n_11223
use :  
dir : i
shape : 
(276450,0):(276550,510) : 1
n_11264
use :  
dir : i
shape : 
(352090,89950):(352600,90050) : 2
n_12153
use :  
dir : i
shape : 
(278650,0):(278750,510) : 1
n_1252
use :  
dir : i
shape : 
(352090,89750):(352600,89850) : 2
n_12825
use :  
dir : i
shape : 
(352090,89550):(352600,89650) : 2
n_1340
use :  
dir : i
shape : 
(352090,89350):(352600,89450) : 2
n_1342
use :  
dir : i
shape : 
(352090,89150):(352600,89250) : 2
n_1354
use :  
dir : i
shape : 
(352090,88950):(352600,89050) : 2
n_15568
use :  
dir : i
shape : 
(258250,0):(258350,510) : 1
n_2401
use :  
dir : i
shape : 
(352090,113150):(352600,113250) : 2
n_8605
use :  
dir : i
shape : 
(251650,159490):(251750,160000) : 1
n_8831
use :  
dir : i
shape : 
(231000,159745):(231200,160000) : 3
n_8832
use :  
dir : i
shape : 
(245050,159490):(245150,160000) : 1
n_8927
use :  
dir : i
shape : 
(231250,0):(231350,510) : 1
n_9116
use :  
dir : i
shape : 
(279050,159490):(279150,160000) : 1
n_9269
use :  
dir : i
shape : 
(165650,0):(165750,510) : 1
n_9372
use :  
dir : i
shape : 
(352090,65950):(352600,66050) : 2
n_9407
use :  
dir : i
shape : 
(92850,0):(92950,510) : 1
n_9586
use :  
dir : i
shape : 
(314850,0):(314950,510) : 1
n_9844
use :  
dir : i
shape : 
(313850,0):(313950,510) : 1
wbu_addr_in_254
use :  
dir : i
shape : 
(303250,159490):(303350,160000) : 1
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__29__Q
use :  
dir : i
shape : 
(133050,0):(133150,510) : 1
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__29__Q
use :  
dir : i
shape : 
(196250,0):(196350,510) : 1
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__27__Q
use :  
dir : i
shape : 
(59250,0):(59350,510) : 1
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__29__Q
use :  
dir : i
shape : 
(258650,0):(258750,510) : 1
h5
--pins(105)
FE_OCPN1988_FE_OFN1264_n_8567
use : z
dir : o
shape : 
(309200,0):(309400,255) : 3
FE_OFN1299_n_8567
use :  
dir : o
shape : 
(117400,0):(117600,255) : 3
FE_OFN1504_n_9531
use :  
dir : o
shape : 
(31850,0):(31950,510) : 1
FE_OFN1675_n_10588
use :  
dir : o
shape : 
(78050,0):(78150,510) : 1
FE_OFN538_n_9895
use : z
dir : o
shape : 
(0,90900):(255,91100) : 2
g57182_da
use : z
dir : o
shape : 
(61650,0):(61750,510) : 1
g57202_db
use : z
dir : o
shape : 
(60850,153490):(60950,154000) : 1
g57368_db
use : z
dir : o
shape : 
(237250,0):(237350,510) : 1
g57569_db
use : Z
dir : o
shape : 
(149450,0):(149550,510) : 1
g57942_sb
use : �
dir : o
shape : 
(71650,0):(71750,510) : 1
g58061_db
use :  
dir : o
shape : 
(74050,153490):(74150,154000) : 1
g58210_db
use : �
dir : o
shape : 
(55050,0):(55150,510) : 1
g58235_db
use : r
dir : o
shape : 
(0,21750):(510,21850) : 2
g58319_db
use :  
dir : o
shape : 
(47850,153490):(47950,154000) : 1
g58425_da
use : �
dir : o
shape : 
(163050,0):(163150,510) : 1
g61860_da
use : �
dir : o
shape : 
(333250,153490):(333350,154000) : 1
n_10554
use :  
dir : o
shape : 
(0,57550):(510,57650) : 2
n_11097
use :  
dir : o
shape : 
(163450,153490):(163550,154000) : 1
n_11198
use :  
dir : o
shape : 
(358490,57150):(359000,57250) : 2
n_11261
use :  
dir : o
shape : 
(358490,57350):(359000,57450) : 2
n_12158
use :  
dir : o
shape : 
(189450,0):(189550,510) : 1
n_12530
use :  
dir : o
shape : 
(109050,153490):(109150,154000) : 1
n_2151
use :  
dir : o
shape : 
(159850,153490):(159950,154000) : 1
n_7842
use :  
dir : o
shape : 
(338250,0):(338350,510) : 1
n_9878
use :  
dir : o
shape : 
(0,57750):(510,57850) : 2
n_9971
use :  
dir : o
shape : 
(256850,0):(256950,510) : 1
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__8__Q
use :  
dir : o
shape : 
(139650,153490):(139750,154000) : 1
pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__22__Q
use :  
dir : o
shape : 
(173650,0):(173750,510) : 1
pci_target_unit_pcit_if_pcir_fifo_data_in_766
use :  
dir : o
shape : 
(136250,153490):(136350,154000) : 1
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__6__Q
use :  
dir : o
shape : 
(216450,0):(216550,510) : 1
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__6__Q
use :  
dir : o
shape : 
(83250,153490):(83350,154000) : 1
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__21__Q
use :  
dir : o
shape : 
(101650,0):(101750,510) : 1
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__6__Q
use :  
dir : o
shape : 
(292050,0):(292150,510) : 1
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__17__Q
use :  
dir : o
shape : 
(129050,0):(129150,510) : 1
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__2__Q
use :  
dir : o
shape : 
(234450,0):(234550,510) : 1
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__6__Q
use :  
dir : o
shape : 
(27450,153490):(27550,154000) : 1
FE_OCPN1987_FE_OFN1264_n_8567
use :  
dir : i
shape : 
(308650,0):(308750,510) : 1
FE_OCP_RBN2065_n_16572
use :  
dir : i
shape : 
(173450,0):(173550,510) : 1
FE_OFN1068_n_8176
use :  
dir : i
shape : 
(358490,90950):(359000,91050) : 2
FE_OFN1077_n_7845
use :  
dir : i
shape : 
(329200,0):(329400,255) : 3
FE_OFN1265_n_8567
use :  
dir : i
shape : 
(358745,57700):(359000,57900) : 2
FE_OFN1271_n_8567
use :  
dir : i
shape : 
(0,90500):(255,90700) : 2
FE_OFN1281_n_8567
use :  
dir : i
shape : 
(64400,0):(64600,255) : 3
FE_OFN1283_n_8567
use :  
dir : i
shape : 
(117650,0):(117750,510) : 1
FE_OFN1322_n_8567
use :  
dir : i
shape : 
(237600,0):(237800,255) : 3
FE_OFN1323_n_8567
use :  
dir : i
shape : 
(274800,0):(275000,255) : 3
FE_OFN1349_n_9163
use :  
dir : i
shape : 
(113850,153490):(113950,154000) : 1
FE_OFN1353_n_15558
use :  
dir : i
shape : 
(147850,0):(147950,510) : 1
FE_OFN1365_n_15587
use :  
dir : i
shape : 
(257450,0):(257550,510) : 1
FE_OFN1376_n_10853
use :  
dir : i
shape : 
(0,57350):(510,57450) : 2
FE_OFN1502_n_9531
use :  
dir : i
shape : 
(32050,0):(32150,510) : 1
FE_OFN1503_n_9531
use :  
dir : i
shape : 
(301450,153490):(301550,154000) : 1
FE_OFN1543_n_9502
use :  
dir : i
shape : 
(358745,126900):(359000,127100) : 2
FE_OFN1544_n_9502
use :  
dir : i
shape : 
(49200,153745):(49400,154000) : 3
FE_OFN1678_n_10588
use :  
dir : i
shape : 
(0,57150):(510,57250) : 2
FE_OFN1682_n_16891
use :  
dir : i
shape : 
(258050,0):(258150,510) : 1
FE_OFN1717_n_16637
use :  
dir : i
shape : 
(113250,153490):(113350,154000) : 1
FE_OFN1842_n_9828
use :  
dir : i
shape : 
(301200,153745):(301400,154000) : 3
FE_OFN222_n_9844
use :  
dir : i
shape : 
(48050,153490):(48150,154000) : 1
FE_OFN239_n_9118
use :  
dir : i
shape : 
(211200,153745):(211400,154000) : 3
FE_OFN521_n_9690
use :  
dir : i
shape : 
(0,21300):(255,21500) : 2
FE_OFN535_n_9895
use :  
dir : i
shape : 
(0,91750):(510,91850) : 2
FE_OFN536_n_9895
use :  
dir : i
shape : 
(88050,0):(88150,510) : 1
FE_OFN551_n_9902
use :  
dir : i
shape : 
(209200,0):(209400,255) : 3
FE_OFN568_n_9694
use :  
dir : i
shape : 
(55400,0):(55600,255) : 3
FE_OFN579_n_9904
use :  
dir : i
shape : 
(74450,153490):(74550,154000) : 1
FE_OFN680_n_8060
use :  
dir : i
shape : 
(238400,153745):(238600,154000) : 3
g57065_db
use :  
dir : i
shape : 
(0,91550):(510,91650) : 2
g57353_da
use :  
dir : i
shape : 
(82250,0):(82350,510) : 1
g57473_db
use :  
dir : i
shape : 
(358490,56950):(359000,57050) : 2
g57932_da
use :  
dir : i
shape : 
(0,56950):(510,57050) : 2
g57942_da
use :  
dir : i
shape : 
(0,91350):(510,91450) : 2
g58425_sb
use :  
dir : i
shape : 
(163450,0):(163550,510) : 1
g61866_da
use :  
dir : i
shape : 
(107650,0):(107750,510) : 1
g62004_sb
use :  
dir : i
shape : 
(292050,153490):(292150,154000) : 1
g62027_db
use :  
dir : i
shape : 
(338650,0):(338750,510) : 1
g65976_da
use :  
dir : i
shape : 
(318050,0):(318150,510) : 1
g65976_db
use :  
dir : i
shape : 
(318250,0):(318350,510) : 1
ispd_clk
use :  
dir : i
shape : 
(102000,0):(102200,255) : 3
n_10151
use :  
dir : i
shape : 
(190250,0):(190350,510) : 1
n_10154
use :  
dir : i
shape : 
(190050,0):(190150,510) : 1
n_10381
use :  
dir : i
shape : 
(291050,0):(291150,510) : 1
n_10414
use :  
dir : i
shape : 
(217450,0):(217550,510) : 1
n_10426
use :  
dir : i
shape : 
(28450,153490):(28550,154000) : 1
n_10588
use :  
dir : i
shape : 
(78250,0):(78350,510) : 1
n_11040
use :  
dir : i
shape : 
(110650,153490):(110750,154000) : 1
n_11041
use :  
dir : i
shape : 
(110050,153490):(110150,154000) : 1
n_11572
use :  
dir : i
shape : 
(130050,0):(130150,510) : 1
n_11773
use :  
dir : i
shape : 
(109650,153490):(109750,154000) : 1
n_12548
use :  
dir : i
shape : 
(137250,153490):(137350,154000) : 1
n_1851
use :  
dir : i
shape : 
(333450,153490):(333550,154000) : 1
n_2053
use :  
dir : i
shape : 
(189200,153745):(189400,154000) : 3
n_2299
use :  
dir : i
shape : 
(173200,153745):(173400,154000) : 3
n_7853
use :  
dir : i
shape : 
(140650,153490):(140750,154000) : 1
n_8407
use :  
dir : i
shape : 
(129200,0):(129400,255) : 3
n_9307
use :  
dir : i
shape : 
(189650,0):(189750,510) : 1
n_9744
use :  
dir : i
shape : 
(61850,0):(61950,510) : 1
pci_target_unit_fifos_pcir_data_in_165
use :  
dir : i
shape : 
(173050,153490):(173150,154000) : 1
pci_target_unit_fifos_pcir_data_in_179
use :  
dir : i
shape : 
(269250,153490):(269350,154000) : 1
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__26__Q
use :  
dir : i
shape : 
(41850,0):(41950,510) : 1
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__3__Q
use :  
dir : i
shape : 
(314250,153490):(314350,154000) : 1
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__3__Q
use :  
dir : i
shape : 
(266250,0):(266350,510) : 1
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__3__Q
use :  
dir : i
shape : 
(74250,153490):(74350,154000) : 1
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__17__Q
use :  
dir : i
shape : 
(163250,0):(163350,510) : 1
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__16__Q
use :  
dir : i
shape : 
(0,20950):(510,21050) : 2
h3
--pins(120)
FE_OFN1630_n_9862
use : a
dir : o
shape : 
(85850,177490):(85950,178000) : 1
FE_OFN199_n_9228
use :  
dir : o
shape : 
(0,46500):(255,46700) : 2
FE_RN_189_0
use :  
dir : o
shape : 
(100250,0):(100350,510) : 1
g57181_sb
use :  
dir : o
shape : 
(34850,0):(34950,510) : 1
g57242_db
use :  
dir : o
shape : 
(173450,0):(173550,510) : 1
g57370_da
use :  
dir : o
shape : 
(81650,0):(81750,510) : 1
g57404_db
use :  
dir : o
shape : 
(175050,177490):(175150,178000) : 1
g57508_sb
use :  
dir : o
shape : 
(95050,0):(95150,510) : 1
g57581_db
use :  
dir : o
shape : 
(123850,0):(123950,510) : 1
g57909_da
use :  
dir : o
shape : 
(0,15350):(510,15450) : 2
g57912_db
use :  
dir : o
shape : 
(222850,0):(222950,510) : 1
g58049_da
use :  
dir : o
shape : 
(0,45950):(510,46050) : 2
g58066_da
use :  
dir : o
shape : 
(0,74950):(510,75050) : 2
g58066_db
use :  
dir : o
shape : 
(277850,0):(277950,510) : 1
g58107_da
use :  
dir : o
shape : 
(75650,177490):(75750,178000) : 1
g58339_da
use :  
dir : o
shape : 
(227850,177490):(227950,178000) : 1
g58434_da
use :  
dir : o
shape : 
(134650,0):(134750,510) : 1
g58437_da
use :  
dir : o
shape : 
(184850,0):(184950,510) : 1
n_10060
use :  
dir : o
shape : 
(161050,0):(161150,510) : 1
n_10608
use :  
dir : o
shape : 
(121250,0):(121350,510) : 1
n_11362
use :  
dir : o
shape : 
(255450,0):(255550,510) : 1
n_11544
use :  
dir : o
shape : 
(250250,0):(250350,510) : 1
n_11582
use :  
dir : o
shape : 
(276250,0):(276350,510) : 1
n_12129
use :  
dir : o
shape : 
(75050,0):(75150,510) : 1
n_12140
use :  
dir : o
shape : 
(21050,0):(21150,510) : 1
n_9427
use :  
dir : o
shape : 
(116850,177490):(116950,178000) : 1
n_9435
use :  
dir : o
shape : 
(64250,177490):(64350,178000) : 1
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__35__Q
use :  
dir : o
shape : 
(0,102950):(510,103050) : 2
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__8__Q
use :  
dir : o
shape : 
(233850,177490):(233950,178000) : 1
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__0__Q
use :  
dir : o
shape : 
(313050,0):(313150,510) : 1
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__33__Q
use :  
dir : o
shape : 
(171250,177490):(171350,178000) : 1
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__35__Q
use :  
dir : o
shape : 
(45450,177490):(45550,178000) : 1
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__14__Q
use :  
dir : o
shape : 
(150250,177490):(150350,178000) : 1
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__32__Q
use :  
dir : o
shape : 
(202850,0):(202950,510) : 1
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__20__Q
use :  
dir : o
shape : 
(100050,177490):(100150,178000) : 1
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__35__Q
use :  
dir : o
shape : 
(56050,0):(56150,510) : 1
wishbone_slave_unit_pcim_if_wbw_addr_data_in_393
use :  
dir : o
shape : 
(107050,0):(107150,510) : 1
wishbone_slave_unit_pcim_if_wbw_addr_data_in_397
use :  
dir : o
shape : 
(0,133150):(510,133250) : 2
wishbone_slave_unit_pcim_if_wbw_addr_data_in_398
use :  
dir : o
shape : 
(0,163150):(510,163250) : 2
wishbone_slave_unit_pcim_if_wbw_addr_data_in_403
use :  
dir : o
shape : 
(0,46150):(510,46250) : 2
FE_OCPN1936_n_15566
use :  
dir : i
shape : 
(57200,0):(57400,255) : 3
FE_OCP_RBN2062_n_16572
use :  
dir : i
shape : 
(98450,0):(98550,510) : 1
FE_OFN1257_n_8567
use :  
dir : i
shape : 
(271000,0):(271200,255) : 3
FE_OFN1273_n_8567
use :  
dir : i
shape : 
(0,73900):(255,74100) : 2
FE_OFN1274_n_8567
use :  
dir : i
shape : 
(356145,102900):(356400,103100) : 2
FE_OFN1285_n_8567
use :  
dir : i
shape : 
(0,74300):(255,74500) : 2
FE_OFN1286_n_8567
use :  
dir : i
shape : 
(144200,177745):(144400,178000) : 3
FE_OFN1288_n_8567
use :  
dir : i
shape : 
(163800,177745):(164000,178000) : 3
FE_OFN1289_n_8567
use :  
dir : i
shape : 
(35000,0):(35200,255) : 3
FE_OFN1292_n_8567
use :  
dir : i
shape : 
(95200,0):(95400,255) : 3
FE_OFN1308_n_8567
use :  
dir : i
shape : 
(0,7500):(255,7700) : 2
FE_OFN1311_n_8567
use :  
dir : i
shape : 
(231000,0):(231200,255) : 3
FE_OFN1312_n_8567
use :  
dir : i
shape : 
(356145,132900):(356400,133100) : 2
FE_OFN1319_n_8567
use :  
dir : i
shape : 
(124200,0):(124400,255) : 3
FE_OFN1320_n_8567
use :  
dir : i
shape : 
(238400,177745):(238600,178000) : 3
FE_OFN1354_n_15558
use :  
dir : i
shape : 
(122050,0):(122150,510) : 1
FE_OFN1355_n_15558
use :  
dir : i
shape : 
(99050,0):(99150,510) : 1
FE_OFN1367_n_15587
use :  
dir : i
shape : 
(85050,0):(85150,510) : 1
FE_OFN1368_n_15587
use :  
dir : i
shape : 
(63450,0):(63550,510) : 1
FE_OFN1378_n_10853
use :  
dir : i
shape : 
(207650,0):(207750,510) : 1
FE_OFN1505_n_9531
use :  
dir : i
shape : 
(25250,177490):(25350,178000) : 1
FE_OFN1537_n_9428
use :  
dir : i
shape : 
(105650,0):(105750,510) : 1
FE_OFN1538_n_9428
use :  
dir : i
shape : 
(183000,0):(183200,255) : 3
FE_OFN1565_n_9477
use :  
dir : i
shape : 
(356145,44900):(356400,45100) : 2
FE_OFN1629_n_9862
use :  
dir : i
shape : 
(86050,177490):(86150,178000) : 1
FE_OFN1677_n_10588
use :  
dir : i
shape : 
(207050,0):(207150,510) : 1
FE_OFN1685_n_16891
use :  
dir : i
shape : 
(85650,0):(85750,510) : 1
FE_OFN1688_n_15534
use :  
dir : i
shape : 
(210050,177490):(210150,178000) : 1
FE_OFN1693_n_16992
use :  
dir : i
shape : 
(210650,177490):(210750,178000) : 1
FE_OFN198_n_9228
use :  
dir : i
shape : 
(0,45750):(510,45850) : 2
FE_OFN201_n_9140
use :  
dir : i
shape : 
(263000,177745):(263200,178000) : 3
FE_OFN203_n_9865
use :  
dir : i
shape : 
(356145,45300):(356400,45500) : 2
FE_OFN210_n_9858
use :  
dir : i
shape : 
(239250,0):(239350,510) : 1
FE_OFN212_n_9124
use :  
dir : i
shape : 
(145400,0):(145600,255) : 3
FE_OFN216_n_9889
use :  
dir : i
shape : 
(0,14900):(255,15100) : 2
FE_OFN254_n_9868
use :  
dir : i
shape : 
(82000,177745):(82200,178000) : 3
FE_OFN268_n_9884
use :  
dir : i
shape : 
(0,45300):(255,45500) : 2
FE_OFN539_n_9895
use :  
dir : i
shape : 
(356145,74700):(356400,74900) : 2
FE_OFN548_n_9502
use :  
dir : i
shape : 
(219200,0):(219400,255) : 3
FE_OFN554_n_9902
use :  
dir : i
shape : 
(231400,0):(231600,255) : 3
FE_OFN560_n_9531
use :  
dir : i
shape : 
(82400,177745):(82600,178000) : 3
FE_OFN571_n_9694
use :  
dir : i
shape : 
(0,15700):(255,15900) : 2
FE_OFN572_n_9694
use :  
dir : i
shape : 
(274800,177745):(275000,178000) : 3
FE_OFN576_n_9687
use :  
dir : i
shape : 
(0,103300):(255,103500) : 2
FE_OFN580_n_9904
use :  
dir : i
shape : 
(278200,0):(278400,255) : 3
FE_OFN581_n_9904
use :  
dir : i
shape : 
(75200,0):(75400,255) : 3
g57213_db
use :  
dir : i
shape : 
(250650,0):(250750,510) : 1
g57221_da
use :  
dir : i
shape : 
(119050,177490):(119150,178000) : 1
g57544_da
use :  
dir : i
shape : 
(55450,177490):(55550,178000) : 1
g57944_da
use :  
dir : i
shape : 
(355890,103350):(356400,103450) : 2
g58060_da
use :  
dir : i
shape : 
(124450,0):(124550,510) : 1
g58073_db
use :  
dir : i
shape : 
(237250,0):(237350,510) : 1
g58333_da
use :  
dir : i
shape : 
(77650,177490):(77750,178000) : 1
g58333_db
use :  
dir : i
shape : 
(77850,177490):(77950,178000) : 1
g58341_sb
use :  
dir : i
shape : 
(330450,0):(330550,510) : 1
g58402_db
use :  
dir : i
shape : 
(64650,177490):(64750,178000) : 1
g58438_db
use :  
dir : i
shape : 
(201050,0):(201150,510) : 1
ispd_clk
use :  
dir : i
shape : 
(0,46900):(255,47100) : 2
n_10002
use :  
dir : i
shape : 
(21650,0):(21750,510) : 1
n_11259
use :  
dir : i
shape : 
(234850,177490):(234950,178000) : 1
n_11337
use :  
dir : i
shape : 
(162850,177490):(162950,178000) : 1
n_11516
use :  
dir : i
shape : 
(186250,177490):(186350,178000) : 1
n_12841
use :  
dir : i
shape : 
(0,44950):(510,45050) : 2
n_12847
use :  
dir : i
shape : 
(0,162950):(510,163050) : 2
n_12848
use :  
dir : i
shape : 
(0,132950):(510,133050) : 2
n_12852
use :  
dir : i
shape : 
(108050,0):(108150,510) : 1
n_16840
use :  
dir : i
shape : 
(21250,0):(21350,510) : 1
n_16841
use :  
dir : i
shape : 
(22250,0):(22350,510) : 1
n_9551
use :  
dir : i
shape : 
(245250,0):(245350,510) : 1
n_9726
use :  
dir : i
shape : 
(259850,0):(259950,510) : 1
n_9868
use :  
dir : i
shape : 
(182850,0):(182950,510) : 1
n_9908
use :  
dir : i
shape : 
(0,74750):(510,74850) : 2
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__34__Q
use :  
dir : i
shape : 
(63650,0):(63750,510) : 1
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__8__Q
use :  
dir : i
shape : 
(86050,0):(86150,510) : 1
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__8__Q
use :  
dir : i
shape : 
(42650,0):(42750,510) : 1
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__0__Q
use :  
dir : i
shape : 
(297450,0):(297550,510) : 1
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__28__Q
use :  
dir : i
shape : 
(162250,0):(162350,510) : 1
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__10__Q
use :  
dir : i
shape : 
(113450,0):(113550,510) : 1
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__28__Q
use :  
dir : i
shape : 
(134850,0):(134950,510) : 1
wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__1__Q
use :  
dir : i
shape : 
(265850,0):(265950,510) : 1
h2
--pins(154)
FE_OCP_RBN2122_n_16966
use :  
dir : o
shape : 
(0,15550):(510,15650) : 2
FE_OFN741_n_2678
use :  
dir : o
shape : 
(225850,0):(225950,510) : 1
FE_OFN752_n_2547
use :  
dir : o
shape : 
(55650,0):(55750,510) : 1
FE_RN_232_0
use :  
dir : o
shape : 
(360090,162750):(360600,162850) : 2
configuration_pci_err_addr_471
use :  
dir : o
shape : 
(139650,0):(139750,510) : 1
configuration_sync_cache_lsize_to_wb_bits_reg_3__Q
use :  
dir : o
shape : 
(360090,45150):(360600,45250) : 2
g53255_p
use :  
dir : o
shape : 
(46650,0):(46750,510) : 1
g53301_p
use :  
dir : o
shape : 
(110850,177490):(110950,178000) : 1
g61965_da
use :  
dir : o
shape : 
(0,162550):(510,162650) : 2
g62827_da
use :  
dir : o
shape : 
(56650,177490):(56750,178000) : 1
g62837_da
use :  
dir : o
shape : 
(0,132950):(510,133050) : 2
g62837_db
use :  
dir : o
shape : 
(0,133150):(510,133250) : 2
g63077_da
use :  
dir : o
shape : 
(87850,0):(87950,510) : 1
g63080_db
use :  
dir : o
shape : 
(0,72550):(510,72650) : 2
g63568_db
use :  
dir : o
shape : 
(37650,177490):(37750,178000) : 1
g64259_db
use :  
dir : o
shape : 
(0,45150):(510,45250) : 2
g64259_sb
use :  
dir : o
shape : 
(0,103350):(510,103450) : 2
g64301_db
use :  
dir : o
shape : 
(61050,177490):(61150,178000) : 1
g64332_db
use :  
dir : o
shape : 
(0,42950):(510,43050) : 2
g64332_sb
use :  
dir : o
shape : 
(0,45350):(510,45450) : 2
g65212_da
use :  
dir : o
shape : 
(293650,0):(293750,510) : 1
g65234_sb
use :  
dir : o
shape : 
(216850,0):(216950,510) : 1
g65240_db
use :  
dir : o
shape : 
(181650,0):(181750,510) : 1
g66184_p
use :  
dir : o
shape : 
(360090,103950):(360600,104050) : 2
g66726_p
use :  
dir : o
shape : 
(360090,14950):(360600,15050) : 2
n_10825
use :  
dir : o
shape : 
(220250,0):(220350,510) : 1
n_1159
use :  
dir : o
shape : 
(260250,0):(260350,510) : 1
n_1196
use :  
dir : o
shape : 
(360090,102950):(360600,103050) : 2
n_13304
use :  
dir : o
shape : 
(114050,0):(114150,510) : 1
n_13701
use :  
dir : o
shape : 
(31650,0):(31750,510) : 1
n_13859
use :  
dir : o
shape : 
(70050,0):(70150,510) : 1
n_13980
use :  
dir : o
shape : 
(98450,177490):(98550,178000) : 1
n_14413
use :  
dir : o
shape : 
(85850,177490):(85950,178000) : 1
n_14690
use :  
dir : o
shape : 
(162250,177490):(162350,178000) : 1
n_14804
use :  
dir : o
shape : 
(143250,177490):(143350,178000) : 1
n_1507
use :  
dir : o
shape : 
(176450,177490):(176550,178000) : 1
n_1552
use :  
dir : o
shape : 
(360090,104150):(360600,104250) : 2
n_15611
use :  
dir : o
shape : 
(252050,0):(252150,510) : 1
n_16275
use :  
dir : o
shape : 
(290450,177490):(290550,178000) : 1
n_16280
use :  
dir : o
shape : 
(234450,0):(234550,510) : 1
n_16507
use :  
dir : o
shape : 
(205450,0):(205550,510) : 1
n_16748
use :  
dir : o
shape : 
(108200,0):(108400,255) : 3
n_16975
use :  
dir : o
shape : 
(0,15750):(510,15850) : 2
n_177
use :  
dir : o
shape : 
(284650,0):(284750,510) : 1
n_2597
use :  
dir : o
shape : 
(206650,0):(206750,510) : 1
n_2598
use :  
dir : o
shape : 
(209450,0):(209550,510) : 1
n_2729
use :  
dir : o
shape : 
(258050,0):(258150,510) : 1
n_2776
use :  
dir : o
shape : 
(125450,0):(125550,510) : 1
n_3123
use :  
dir : o
shape : 
(360090,103350):(360600,103450) : 2
n_3319
use :  
dir : o
shape : 
(214450,0):(214550,510) : 1
n_3320
use :  
dir : o
shape : 
(193650,0):(193750,510) : 1
n_8498
use :  
dir : o
shape : 
(300650,0):(300750,510) : 1
n_8757
use :  
dir : o
shape : 
(147200,0):(147400,255) : 3
n_8759
use :  
dir : o
shape : 
(102650,0):(102750,510) : 1
n_8800
use :  
dir : o
shape : 
(288450,177490):(288550,178000) : 1
n_8879
use :  
dir : o
shape : 
(146850,0):(146950,510) : 1
n_9175
use :  
dir : o
shape : 
(360090,75350):(360600,75450) : 2
pci_target_unit_fifos_pciw_addr_data_in_121
use :  
dir : o
shape : 
(0,103550):(510,103650) : 2
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__35__Q
use :  
dir : o
shape : 
(0,102950):(510,103050) : 2
pci_target_unit_pcit_if_strd_bc_in
use :  
dir : o
shape : 
(270450,177490):(270550,178000) : 1
pci_target_unit_pcit_if_strd_bc_in_718
use :  
dir : o
shape : 
(203050,177490):(203150,178000) : 1
pci_target_unit_pcit_if_strd_bc_in_719
use :  
dir : o
shape : 
(166450,0):(166550,510) : 1
wbm_sel_o_0_
use :  
dir : o
shape : 
(0,68550):(510,68650) : 2
wbm_sel_o_3_
use :  
dir : o
shape : 
(0,103750):(510,103850) : 2
FE_OCP_RBN2123_n_16966
use :  
dir : i
shape : 
(0,15950):(510,16050) : 2
FE_OFN1017_g64577_p
use :  
dir : i
shape : 
(0,72100):(255,72300) : 2
FE_OFN1019_g64577_p
use :  
dir : i
shape : 
(101600,177745):(101800,178000) : 3
FE_OFN1112_n_3476
use :  
dir : i
shape : 
(119800,0):(120000,255) : 3
FE_OFN1463_n_13736
use :  
dir : i
shape : 
(96850,0):(96950,510) : 1
FE_OFN1520_n_4730
use :  
dir : i
shape : 
(66400,177745):(66600,178000) : 3
FE_OFN1776_n_13971
use :  
dir : i
shape : 
(98600,177745):(98800,178000) : 3
FE_OFN189_n_1193
use :  
dir : i
shape : 
(301250,177490):(301350,178000) : 1
FE_OFN747_n_2678
use :  
dir : i
shape : 
(186400,0):(186600,255) : 3
FE_OFN751_n_2547
use :  
dir : i
shape : 
(55850,0):(55950,510) : 1
FE_OFN860_n_4734
use :  
dir : i
shape : 
(0,133700):(255,133900) : 2
FE_OFN959_n_16760
use :  
dir : i
shape : 
(110450,0):(110550,510) : 1
FE_OFN973_n_4727
use :  
dir : i
shape : 
(0,44500):(255,44700) : 2
FE_RN_285_0
use :  
dir : i
shape : 
(234650,0):(234750,510) : 1
FE_RN_286_0
use :  
dir : i
shape : 
(234850,0):(234950,510) : 1
FE_RN_345_0
use :  
dir : i
shape : 
(311650,0):(311750,510) : 1
FE_RN_427_0
use :  
dir : i
shape : 
(119850,177490):(119950,178000) : 1
configuration_meta_cache_lsize_to_wb_bits_926
use :  
dir : i
shape : 
(360090,44950):(360600,45050) : 2
configuration_sync_cache_lsize_to_wb_bits_reg_2__Q
use :  
dir : i
shape : 
(244650,0):(244750,510) : 1
g60615_db
use :  
dir : i
shape : 
(158450,0):(158550,510) : 1
g63564_sb
use :  
dir : i
shape : 
(161450,177490):(161550,178000) : 1
g65215_da
use :  
dir : i
shape : 
(227650,177490):(227750,178000) : 1
g65225_da
use :  
dir : i
shape : 
(220650,177490):(220750,178000) : 1
g65234_da
use :  
dir : i
shape : 
(227250,0):(227350,510) : 1
ispd_clk
use :  
dir : i
shape : 
(140000,0):(140200,255) : 3
n_1219
use :  
dir : i
shape : 
(176650,177490):(176750,178000) : 1
n_1304
use :  
dir : i
shape : 
(360090,133150):(360600,133250) : 2
n_13122
use :  
dir : i
shape : 
(114250,0):(114350,510) : 1
n_13484
use :  
dir : i
shape : 
(134250,0):(134350,510) : 1
n_1366
use :  
dir : i
shape : 
(360090,103150):(360600,103250) : 2
n_13919
use :  
dir : i
shape : 
(322050,177490):(322150,178000) : 1
n_13955
use :  
dir : i
shape : 
(46850,0):(46950,510) : 1
n_13971
use :  
dir : i
shape : 
(123250,177490):(123350,178000) : 1
n_1435
use :  
dir : i
shape : 
(360090,75150):(360600,75250) : 2
n_14529
use :  
dir : i
shape : 
(301050,177490):(301150,178000) : 1
n_14829
use :  
dir : i
shape : 
(134050,0):(134150,510) : 1
n_14837
use :  
dir : i
shape : 
(102850,0):(102950,510) : 1
n_14895
use :  
dir : i
shape : 
(133650,0):(133750,510) : 1
n_14897
use :  
dir : i
shape : 
(0,72750):(510,72850) : 2
n_15114
use :  
dir : i
shape : 
(32250,0):(32350,510) : 1
n_1513
use :  
dir : i
shape : 
(279450,0):(279550,510) : 1
n_15292
use :  
dir : i
shape : 
(323450,0):(323550,510) : 1
n_15302
use :  
dir : i
shape : 
(258450,0):(258550,510) : 1
n_1551
use :  
dir : i
shape : 
(360090,103750):(360600,103850) : 2
n_15607
use :  
dir : i
shape : 
(278850,0):(278950,510) : 1
n_16205
use :  
dir : i
shape : 
(32450,0):(32550,510) : 1
n_16331
use :  
dir : i
shape : 
(360090,103550):(360600,103650) : 2
n_16738
use :  
dir : i
shape : 
(108450,0):(108550,510) : 1
n_16966
use :  
dir : i
shape : 
(0,15350):(510,15450) : 2
n_16970
use :  
dir : i
shape : 
(0,15150):(510,15250) : 2
n_16974
use :  
dir : i
shape : 
(0,14950):(510,15050) : 2
n_2031
use :  
dir : i
shape : 
(258250,0):(258350,510) : 1
n_2301
use :  
dir : i
shape : 
(360345,74100):(360600,74300) : 2
n_2337
use :  
dir : i
shape : 
(302850,0):(302950,510) : 1
n_2353
use :  
dir : i
shape : 
(297850,0):(297950,510) : 1
n_2599
use :  
dir : i
shape : 
(176650,0):(176750,510) : 1
n_2675
use :  
dir : i
shape : 
(293850,0):(293950,510) : 1
n_2677
use :  
dir : i
shape : 
(167450,0):(167550,510) : 1
n_2678
use :  
dir : i
shape : 
(268650,0):(268750,510) : 1
n_2730
use :  
dir : i
shape : 
(125650,0):(125750,510) : 1
n_2779
use :  
dir : i
shape : 
(360090,74950):(360600,75050) : 2
n_4592
use :  
dir : i
shape : 
(0,162750):(510,162850) : 2
n_5092
use :  
dir : i
shape : 
(0,103150):(510,103250) : 2
n_657
use :  
dir : i
shape : 
(341850,0):(341950,510) : 1
n_7698
use :  
dir : i
shape : 
(360090,132950):(360600,133050) : 2
n_8487
use :  
dir : i
shape : 
(332850,0):(332950,510) : 1
n_8538
use :  
dir : i
shape : 
(298250,0):(298350,510) : 1
n_8819
use :  
dir : i
shape : 
(279250,0):(279350,510) : 1
n_9178
use :  
dir : i
shape : 
(318850,177490):(318950,178000) : 1
output_backup_trdy_out_reg_Q
use :  
dir : i
shape : 
(192650,0):(192750,510) : 1
parchk_pci_ad_reg_in
use :  
dir : i
shape : 
(263650,177490):(263750,178000) : 1
parchk_pci_ad_reg_in_1205
use :  
dir : i
shape : 
(243450,0):(243550,510) : 1
pci_target_unit_del_sync_bc_in
use :  
dir : i
shape : 
(233250,177490):(233350,178000) : 1
pci_target_unit_del_sync_be_out_reg_3__Q
use :  
dir : i
shape : 
(181850,0):(181950,510) : 1
pci_target_unit_fifos_pciw_addr_data_in_123
use :  
dir : i
shape : 
(61250,177490):(61350,178000) : 1
pci_target_unit_fifos_pciw_addr_data_in_126
use :  
dir : i
shape : 
(0,44950):(510,45050) : 2
pci_target_unit_fifos_pciw_cbe_in
use :  
dir : i
shape : 
(0,43150):(510,43250) : 2
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__1__Q
use :  
dir : i
shape : 
(70450,0):(70550,510) : 1
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__32__Q
use :  
dir : i
shape : 
(56850,0):(56950,510) : 1
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__3__Q
use :  
dir : i
shape : 
(83450,0):(83550,510) : 1
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__6__Q
use :  
dir : i
shape : 
(96650,0):(96750,510) : 1
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__32__Q
use :  
dir : i
shape : 
(0,133350):(510,133450) : 2
pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__3__Q
use :  
dir : i
shape : 
(75650,177490):(75750,178000) : 1
pci_target_unit_pcit_if_req_req_pending_in
use :  
dir : i
shape : 
(341650,0):(341750,510) : 1
pci_target_unit_pcit_if_strd_bc_in_717
use :  
dir : i
shape : 
(290250,177490):(290350,178000) : 1
pci_target_unit_wbm_sm_pciw_fifo_addr_data_in
use :  
dir : i
shape : 
(124650,177490):(124750,178000) : 1
pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_50
use :  
dir : i
shape : 
(163450,177490):(163550,178000) : 1
pciu_cache_lsize_not_zero_in
use :  
dir : i
shape : 
(205850,0):(205950,510) : 1
wbm_adr_o_0_
use :  
dir : i
shape : 
(92450,0):(92550,510) : 1
wbm_adr_o_1_
use :  
dir : i
shape : 
(0,122550):(510,122650) : 2
ms00f80
--pins(3)
o
use :  
dir : o
shape : 
(50,500):(150,1500) : 1
ck
use :  
dir : i
shape : 
(450,500):(550,1500) : 0
d
use :  
dir : i
shape : 
(1050,500):(1150,1500) : 0
in01f01
--pins(2)
o
use :  
dir : o
shape : 
(50,500):(150,1500) : 0
a
use :  
dir : i
shape : 
(250,500):(350,1500) : 0
no02f01
--pins(3)
o
use :  
dir : o
shape : 
(50,500):(150,1500) : 0
a
use :  
dir : i
shape : 
(250,500):(350,1500) : 0
b
use : z
dir : i
shape : 
(450,500):(550,1500) : 0
na02f01
--pins(3)
o
use :  
dir : o
shape : 
(50,500):(150,1500) : 0
a
use :  
dir : i
shape : 
(250,500):(350,1500) : 0
b
use :  
dir : i
shape : 
(450,500):(550,1500) : 0
ao12f01
--pins(4)
o
use :  
dir : o
shape : 
(50,500):(150,1500) : 0
a
use :  
dir : i
shape : 
(250,500):(350,1500) : 0
b
use : 
dir : i
shape : 
(650,500):(750,1500) : 0
c
use : �
dir : i
shape : 
(850,500):(950,1500) : 0
na03f01
--pins(4)
o
use :  
dir : o
shape : 
(50,500):(150,1500) : 0
a
use :  
dir : i
shape : 
(250,500):(350,1500) : 0
b
use :  
dir : i
shape : 
(650,500):(750,1500) : 0
c
use :  
dir : i
shape : 
(850,500):(950,1500) : 0
oa12f01
--pins(4)
o
use :  
dir : o
shape : 
(50,500):(150,1500) : 0
a
use :  
dir : i
shape : 
(250,500):(350,1500) : 0
b
use :  
dir : i
shape : 
(650,500):(750,1500) : 0
c
use :  
dir : i
shape : 
(850,500):(950,1500) : 0
na04m01
--pins(5)
o
use :  
dir : o
shape : 
(50,500):(150,1500) : 0
a
use :  
dir : i
shape : 
(250,500):(350,1500) : 0
b
use :  
dir : i
shape : 
(650,500):(750,1500) : 0
c
use :  
dir : i
shape : 
(850,500):(950,1500) : 0
d
use :  
dir : i
shape : 
(1250,500):(1350,1500) : 0
no04s01
--pins(5)
o
use :  
dir : o
shape : 
(50,500):(150,1500) : 0
a
use :  
dir : i
shape : 
(250,500):(350,1500) : 0
b
use :  
dir : i
shape : 
(650,500):(750,1500) : 0
c
use :  
dir : i
shape : 
(850,500):(950,1500) : 0
d
use :  
dir : i
shape : 
(1250,500):(1350,1500) : 0
no03m01
--pins(4)
o
use :  
dir : o
shape : 
(50,500):(150,1500) : 0
a
use :  
dir : i
shape : 
(250,500):(350,1500) : 0
b
use :  
dir : i
shape : 
(650,500):(750,1500) : 0
c
use :  
dir : i
shape : 
(850,500):(950,1500) : 0
ao22s01
--pins(5)
o
use :  
dir : o
shape : 
(50,500):(150,1500) : 0
a
use :  
dir : i
shape : 
(250,500):(350,1500) : 0
b
use :  
dir : i
shape : 
(650,500):(750,1500) : 0
c
use :  
dir : i
shape : 
(850,500):(950,1500) : 0
d
use :  
dir : i
shape : 
(1250,500):(1350,1500) : 0
oa22f01
--pins(5)
o
use :  
dir : o
shape : 
(1350,950):(1550,1050) : 1
(1250,500):(1350,1050) : 1
a
use :  
dir : i
shape : 
(250,500):(350,1500) : 0
b
use :  
dir : i
shape : 
(650,500):(750,1500) : 0
c
use :  
dir : i
shape : 
(850,500):(950,1500) : 0
d
use :  
dir : i
shape : 
(50,500):(150,1500) : 0
metal1 (H) p200,200 w100 s110 a41000 prefer: srt200 stp200 num4529 wrong: srt100 stp200 num4530
metal2 (V) p200,200 w100 s120 a51000 prefer: srt100 stp200 num4530 wrong: srt200 stp200 num4529
metal3 (H) p200,200 w100 s120 a51000 prefer: srt200 stp200 num4529 wrong: srt100 stp200 num4530
metal4 (V) p200,200 w100 s120 a51000 prefer: srt100 stp200 num4530 wrong: srt200 stp200 num4529
metal5 (H) p200,200 w100 s120 a51000 prefer: srt200 stp200 num4529 wrong: srt100 stp200 num4530
