net1237
net1240
net1233
net1236
net1234
net1232
net1231
net1239
net1235
net1238
net1230
AOI221X2
--pins(8)
A0
use : s
dir : i
shape : 
(470,1250):(730,1430) : 0
(570,1220):(1920,1380) : 0
(570,1220):(730,1430) : 0
(470,1250):(1920,1380) : 0
A1
use : s
dir : i
shape : 
(1320,1530):(1480,2130) : 0
B0
use : s
dir : i
shape : 
(3270,1250):(3530,1430) : 0
(2480,1270):(3870,1430) : 0
B1
use : s
dir : i
shape : 
(2870,1630):(3870,1790) : 0
C0
use : s
dir : i
shape : 
(4130,1630):(5130,1790) : 0
VDD
use : p
dir : b
shape : 
(0,3300):(5200,3420) : 0
VSS
use : g
dir : b
shape : 
(0,0):(5200,120) : 0
Y
use : s
dir : o
shape : 
(2120,1580):(2280,1840) : 0
(4440,1990):(4560,2270) : 0
(2160,1990):(4560,2110) : 0
(2160,900):(2280,2110) : 0
(1210,900):(4340,1020) : 0
NAND3X2
--pins(6)
A
use : s
dir : i
shape : 
(520,1200):(740,1470) : 0
(2480,990):(2600,1470) : 0
(620,990):(2600,1110) : 0
(620,990):(740,1470) : 0
B
use : s
dir : i
shape : 
(2120,1310):(2280,1840) : 0
(940,1310):(2280,1430) : 0
C
use : s
dir : i
shape : 
(1040,1630):(1530,1910) : 0
(1040,1630):(1920,1790) : 0
VDD
use : p
dir : b
shape : 
(0,3300):(3200,3420) : 0
VSS
use : g
dir : b
shape : 
(0,0):(3200,120) : 0
Y
use : s
dir : o
shape : 
(2870,2010):(3130,2230) : 0
(720,2110):(860,2670) : 0
(3010,670):(3130,2230) : 0
(2380,2110):(2500,2670) : 0
(1590,670):(3130,790) : 0
(1560,2110):(1680,2670) : 0
(720,2110):(3130,2230) : 0
AOI222X1
--pins(9)
A0
use : s
dir : i
shape : 
(520,980):(680,1980) : 0
A1
use : s
dir : i
shape : 
(920,440):(1090,1430) : 0
B0
use : s
dir : i
shape : 
(1760,1720):(2190,2200) : 0
(1720,1510):(1880,1840) : 0
(1760,1510):(1880,2200) : 0
(1720,1720):(2190,1840) : 0
B1
use : s
dir : i
shape : 
(1320,1240):(1520,1840) : 0
(1360,1240):(1520,2200) : 0
C0
use : s
dir : i
shape : 
(2390,1580):(2680,1840) : 0
(2390,1580):(2550,2450) : 0
C1
use : s
dir : i
shape : 
(2880,1240):(3080,2200) : 0
VDD
use : p
dir : b
shape : 
(0,3300):(3600,3420) : 0
VSS
use : g
dir : b
shape : 
(0,0):(3600,120) : 0
Y
use : s
dir : o
shape : 
(2900,820):(3440,1040) : 0
(3320,1960):(3480,2520) : 0
(3320,820):(3440,2520) : 0
(2750,2400):(3480,2520) : 0
(2750,2400):(2870,2640) : 0
(1520,920):(3440,1040) : 0
(1520,760):(1640,1040) : 0
NOR4X4
--pins(7)
A
use : s
dir : i
shape : 
(1720,1510):(1880,1900) : 0
(700,1740):(1880,1900) : 0
B
use : s
dir : i
shape : 
(3450,1510):(3610,1790) : 0
(2480,1630):(3610,1790) : 0
C
use : s
dir : i
shape : 
(4870,1550):(5140,1790) : 0
(4220,1630):(5140,1790) : 0
D
use : s
dir : i
shape : 
(6210,1550):(6370,1790) : 0
(5670,1630):(6840,1790) : 0
VDD
use : p
dir : b
shape : 
(0,3300):(7600,3420) : 0
VSS
use : g
dir : b
shape : 
(0,0):(7600,120) : 0
Y
use : s
dir : o
shape : 
(2120,1580):(2280,1840) : 0
(6920,1030):(7040,1310) : 0
(6810,1990):(6930,2270) : 0
(6100,1030):(6220,1310) : 0
(5990,1990):(6110,2270) : 0
(5280,1030):(5400,1310) : 0
(4460,1030):(4580,1310) : 0
(3640,1030):(3760,1310) : 0
(2820,1030):(2940,1310) : 0
(2160,1990):(6930,2110) : 0
(2160,1190):(2280,2110) : 0
(2000,1030):(2120,1310) : 0
(1180,1190):(7040,1310) : 0
(1180,1030):(1300,1310) : 0
NOR4X2
--pins(7)
A
use : s
dir : i
shape : 
(3320,1960):(3480,2370) : 0
(3360,1640):(3480,2370) : 0
(520,2250):(3480,2370) : 0
(520,1640):(640,2370) : 0
B
use : s
dir : i
shape : 
(920,1580):(1080,1840) : 0
(2870,1690):(2990,2050) : 0
(960,1930):(2990,2050) : 0
(960,1580):(1080,2050) : 0
(840,1670):(1080,1790) : 0
C
use : s
dir : i
shape : 
(2550,1250):(3130,1410) : 0
(2550,1250):(2670,1730) : 0
(1280,1610):(2670,1730) : 0
D
use : s
dir : i
shape : 
(1280,1250):(2280,1410) : 0
VDD
use : p
dir : b
shape : 
(0,3300):(4000,3420) : 0
VSS
use : g
dir : b
shape : 
(0,0):(4000,120) : 0
Y
use : s
dir : o
shape : 
(3720,2340):(3880,2690) : 0
(3190,890):(3430,1050) : 0
(2310,890):(2550,1050) : 0
(1430,890):(1670,1050) : 0
(3760,930):(3880,2690) : 0
(2020,2570):(3880,2690) : 0
(690,930):(3880,1050) : 0
(550,890):(790,1010) : 0
NAND4X2
--pins(7)
A
use : s
dir : i
shape : 
(3720,1640):(3880,2370) : 0
(520,2250):(3880,2370) : 0
(520,1640):(640,2370) : 0
B
use : s
dir : i
shape : 
(920,1580):(1080,1840) : 0
(3200,1690):(3320,2050) : 0
(960,1930):(3320,2050) : 0
(960,1580):(1080,2050) : 0
(840,1670):(1080,1790) : 0
C
use : s
dir : i
shape : 
(2470,1250):(2790,1410) : 0
(2670,1250):(2790,1730) : 0
(1370,1610):(2790,1730) : 0
D
use : s
dir : i
shape : 
(1720,1250):(2270,1410) : 0
(1720,800):(1880,1410) : 0
VDD
use : p
dir : b
shape : 
(0,3300):(4400,3420) : 0
VSS
use : g
dir : b
shape : 
(0,0):(4400,120) : 0
Y
use : s
dir : o
shape : 
(4120,2340):(4280,2690) : 0
(4120,930):(4240,2690) : 0
(3460,2570):(3580,2810) : 0
(2520,2570):(2640,2810) : 0
(2370,930):(4240,1050) : 0
(2140,890):(2470,1010) : 0
(1580,2570):(1700,2810) : 0
(640,2570):(4280,2690) : 0
(640,2570):(760,2810) : 0
BUFX3
--pins(4)
A
use : s
dir : i
shape : 
(1720,1440):(1880,2440) : 0
VDD
use : p
dir : b
shape : 
(0,3300):(2400,3420) : 0
VSS
use : g
dir : b
shape : 
(0,0):(2400,120) : 0
Y
use : s
dir : o
shape : 
(520,1960):(680,2220) : 0
(1250,2100):(1370,2880) : 0
(1170,690):(1290,930) : 0
(1080,810):(1290,930) : 0
(1080,810):(1200,1240) : 0
(520,1120):(640,2220) : 0
(430,2100):(1370,2220) : 0
(430,2100):(550,2880) : 0
(350,1120):(1200,1240) : 0
(350,960):(470,1240) : 0
AOI22X2
--pins(7)
A0
use : s
dir : i
shape : 
(1680,1270):(2130,1430) : 0
(1680,1150):(1840,1430) : 0
(960,1150):(1840,1310) : 0
(960,1150):(1120,1410) : 0
(470,1250):(1120,1410) : 0
A1
use : s
dir : i
shape : 
(1310,1430):(1490,1920) : 0
B0
use : s
dir : i
shape : 
(3680,1160):(3920,1790) : 0
(3680,1630):(4330,1790) : 0
(3000,1160):(3920,1280) : 0
(3000,1160):(3120,1430) : 0
(2650,1310):(3120,1430) : 0
B1
use : s
dir : i
shape : 
(3320,1480):(3480,2060) : 0
VDD
use : p
dir : b
shape : 
(0,3300):(4400,3420) : 0
VSS
use : g
dir : b
shape : 
(0,0):(4400,120) : 0
Y
use : s
dir : o
shape : 
(2070,1630):(2450,1790) : 0
(3680,1990):(3800,2330) : 0
(2860,2210):(3800,2330) : 0
(2860,1670):(2980,2330) : 0
(2330,830):(2450,1790) : 0
(2070,1670):(2980,1790) : 0
(1420,830):(3370,950) : 0
OR4X1
--pins(7)
A
use : s
dir : i
shape : 
(2120,950):(2280,1530) : 0
(1700,1370):(2280,1530) : 0
B
use : s
dir : i
shape : 
(920,1960):(1180,2140) : 0
(1020,1320):(1180,2140) : 0
(920,1960):(1080,2220) : 0
C
use : s
dir : i
shape : 
(660,1180):(820,1740) : 0
(520,1580):(820,1740) : 0
(520,1580):(680,2040) : 0
D
use : s
dir : i
shape : 
(120,1180):(320,1590) : 0
(60,1470):(240,2080) : 0
(120,1180):(240,2080) : 0
(60,1470):(320,1590) : 0
VDD
use : p
dir : b
shape : 
(0,3300):(2800,3420) : 0
VSS
use : g
dir : b
shape : 
(0,0):(2800,120) : 0
Y
use : s
dir : o
shape : 
(2480,820):(2680,1080) : 0
(2480,790):(2600,2770) : 0
NAND3X1
--pins(6)
A
use : s
dir : i
shape : 
(520,1200):(680,2200) : 0
B
use : s
dir : i
shape : 
(960,960):(1120,1780) : 0
(920,820):(1080,1080) : 0
(960,820):(1080,1780) : 0
(920,960):(1120,1080) : 0
C
use : s
dir : i
shape : 
(1320,1200):(1480,2200) : 0
VDD
use : p
dir : b
shape : 
(0,3300):(2000,3420) : 0
VSS
use : g
dir : b
shape : 
(0,0):(2000,120) : 0
Y
use : s
dir : o
shape : 
(1720,2400):(1880,2980) : 0
(1720,880):(1840,2980) : 0
(1490,880):(1840,1000) : 0
(1490,760):(1610,1000) : 0
(850,2400):(1880,2520) : 0
(850,2400):(970,2960) : 0
NOR2X1
--pins(5)
A
use : s
dir : i
shape : 
(520,1140):(680,2140) : 0
B
use : s
dir : i
shape : 
(920,1960):(1120,2170) : 0
(960,1460):(1120,2170) : 0
(920,1960):(1080,2420) : 0
(960,1460):(1080,2420) : 0
VDD
use : p
dir : b
shape : 
(0,3300):(1600,3420) : 0
VSS
use : g
dir : b
shape : 
(0,0):(1600,120) : 0
Y
use : s
dir : o
shape : 
(1320,1200):(1480,1460) : 0
(1320,1140):(1440,2580) : 0
(920,1140):(1440,1260) : 0
(920,980):(1040,1260) : 0
AOI221X1
--pins(8)
A0
use : s
dir : i
shape : 
(520,900):(680,1900) : 0
A1
use : s
dir : i
shape : 
(920,440):(1080,1440) : 0
B0
use : s
dir : i
shape : 
(2120,1160):(2280,2160) : 0
B1
use : s
dir : i
shape : 
(1720,1160):(1880,2160) : 0
C0
use : s
dir : i
shape : 
(2520,1300):(2760,1460) : 0
(2520,1160):(2680,2080) : 0
VDD
use : p
dir : b
shape : 
(0,3300):(3600,3420) : 0
VSS
use : g
dir : b
shape : 
(0,0):(3600,120) : 0
Y
use : s
dir : o
shape : 
(2920,440):(3080,960) : 0
(2960,440):(3080,2920) : 0
(1740,840):(3080,960) : 0
(1600,800):(1840,920) : 0
NAND4X1
--pins(7)
A
use : s
dir : i
shape : 
(460,1300):(680,1840) : 0
(60,1680):(680,1840) : 0
B
use : s
dir : i
shape : 
(960,920):(1120,1780) : 0
(920,920):(1120,1080) : 0
(920,820):(1080,1080) : 0
(960,820):(1080,1780) : 0
C
use : s
dir : i
shape : 
(1320,440):(1480,1660) : 0
D
use : s
dir : i
shape : 
(1720,820):(1880,1820) : 0
VDD
use : p
dir : b
shape : 
(0,3300):(2400,3420) : 0
VSS
use : g
dir : b
shape : 
(0,0):(2400,120) : 0
Y
use : s
dir : o
shape : 
(2080,1580):(2280,2160) : 0
(2080,1080):(2200,2160) : 0
(1580,2040):(1700,2600) : 0
(740,2040):(2280,2160) : 0
(740,2040):(860,2600) : 0
AOI22X1
--pins(7)
A0
use : s
dir : i
shape : 
(520,1200):(680,2200) : 0
A1
use : s
dir : i
shape : 
(960,540):(1120,1400) : 0
(920,540):(1120,700) : 0
(920,440):(1080,700) : 0
(960,440):(1080,1400) : 0
B0
use : s
dir : i
shape : 
(2120,900):(2280,1900) : 0
B1
use : s
dir : i
shape : 
(1720,820):(1880,1820) : 0
VDD
use : p
dir : b
shape : 
(0,3300):(2800,3420) : 0
VSS
use : g
dir : b
shape : 
(0,0):(2800,120) : 0
Y
use : s
dir : o
shape : 
(1320,1960):(1480,2220) : 0
(1870,2100):(1990,2380) : 0
(1360,740):(1480,2220) : 0
(1320,2100):(1990,2220) : 0
BUFX6
--pins(4)
A
use : s
dir : i
shape : 
(2920,1140):(3080,2140) : 0
VDD
use : p
dir : b
shape : 
(0,3300):(3600,3420) : 0
VSS
use : g
dir : b
shape : 
(0,0):(3600,120) : 0
Y
use : s
dir : o
shape : 
(120,1580):(280,1950) : 0
(120,700):(260,2740) : 0
(1780,1830):(1900,2740) : 0
(1780,700):(1900,1310) : 0
(960,1830):(1080,2740) : 0
(960,700):(1080,1310) : 0
(120,1830):(1900,1950) : 0
(120,1190):(1900,1310) : 0
AO22XL
--pins(7)
A0
use : s
dir : i
shape : 
(520,1200):(680,2200) : 0
A1
use : s
dir : i
shape : 
(920,460):(1080,1460) : 0
B0
use : s
dir : i
shape : 
(2120,1580):(2280,2460) : 0
(2000,1580):(2280,1740) : 0
B1
use : s
dir : i
shape : 
(1320,1190):(1480,2190) : 0
VDD
use : p
dir : b
shape : 
(0,3300):(3200,3420) : 0
VSS
use : g
dir : b
shape : 
(0,0):(3200,120) : 0
Y
use : s
dir : o
shape : 
(2520,1820):(3020,1980) : 0
(2520,1200):(2680,1980) : 0
(2500,1200):(2680,1360) : 0
(2500,810):(2660,1360) : 0
(2520,810):(2660,1980) : 0
Metal1 (H) p380,380 w120 s120 a80000 prefer: srt72010 stp380 num51 wrong: srt83800 stp400 num52
Metal2 (V) p400,400 w140 s140 a80000 prefer: srt83800 stp400 num52 wrong: srt72010 stp380 num51
Metal3 (H) p400,400 w140 s140 a80000 prefer: srt72010 stp380 num51 wrong: srt83800 stp400 num52
Metal4 (V) p400,400 w140 s140 a80000 prefer: srt83800 stp400 num52 wrong: srt72010 stp380 num51
Metal5 (H) p400,400 w140 s140 a80000 prefer: srt72010 stp380 num51 wrong: srt83800 stp400 num52
Metal6 (V) p400,400 w140 s140 a80000 prefer: srt83800 stp400 num52 wrong: srt72010 stp380 num51
Metal7 (H) p400,400 w140 s140 a80000 prefer: srt72580 stp570 num33 wrong: srt83800 stp400 num52
Metal8 (V) p400,400 w140 s140 a80000 prefer: srt83800 stp400 num52 wrong: srt72580 stp570 num33
Metal9 (H) p660,660 w140 s140 a80000 prefer: srt72770 stp760 num25 wrong: srt83800 stp400 num52
