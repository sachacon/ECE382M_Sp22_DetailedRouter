net5719
net5021
net5788
net7311
net5532
net6432
net3162
net3947
net7537
net4683
net6796
net6550
net446
net736
net622
net8634
net405
net2142
net8628
net7628
net8428
net4795
net3583
net4502
net7701
net148
net7772
net7563
net796
net8098
net830
net6107
net6821
net6133
net1530
net929
net1793
net6856
net7438
net7323
net7004
net4239
net4631
net4264
net7968
net4057
net2649
net1658
net2304
net6657
net5382
net2442
net7649
net5074
net6
net7026
net6176
net8952
net8951
net8950
net8949
net8948
net8947
net8946
net8945
net8944
net8943
net8942
net8941
net8940
net8939
net8938
net8937
net8936
net8935
net8934
net8933
net8932
net8931
net8930
net8929
net8928
net8927
net8926
net8925
net8924
net8923
net8922
net8921
net8920
net8919
net8918
net8917
net8916
net8915
net8914
net8913
net8912
net8911
net8910
net8909
net8908
net8907
net8906
net8905
net8904
net8903
net8902
net8901
net8900
net8899
net8898
net8897
net8896
net8895
net8894
net8893
net8892
net8891
net8890
net8889
net8888
net8887
net8886
net8885
net8884
net8883
net8882
net8881
net8880
net8879
net8878
net8877
net8876
net8875
net8874
net8873
net8872
net8871
net8870
net8869
net8868
net8867
net8866
net8865
net8864
net8863
net8862
net8861
net8860
net8859
net8858
net8857
net8856
net8855
net8854
net8853
net8852
net8851
net8850
net8849
net8848
net8847
net8846
net8845
net8844
net8843
net8842
net8841
net8840
net8839
net8838
net8837
net8836
net8835
net8834
net8833
net8832
net8831
net8830
net8829
net8828
net8827
net8826
net8825
net8824
net8823
net8822
net8821
net8820
net8819
net8818
net8817
net8816
net8815
net8814
net8813
net8812
net8811
net8810
net8809
net8808
net8807
net8806
net8805
net8804
net8803
net8802
net8801
net8800
net8799
net8798
net8797
net8796
net8795
net8794
net8793
net8792
net8791
net8790
net8789
net8788
net8787
net8786
net8785
net8784
net8783
net8782
net8781
net8780
net8779
net8778
net8777
net8776
net8775
net8774
net8773
net8772
net8771
net8770
net8769
net8768
net8767
net8766
net8765
net8764
net8763
net8762
net8761
net8760
net8759
net8758
net8757
net8756
net8755
net8754
net8753
net8752
net8751
net8750
net8749
net8748
net8747
net8746
net8745
net8744
net8743
net8742
net8741
net8740
net8739
net8738
net8737
net8736
net8735
net8734
net8733
net8732
net8731
net8730
net8729
net8728
net8727
net8726
net8725
net8724
net8723
net8722
net8721
net8720
net8719
net8718
net8717
net8716
net8715
net8714
net8713
net8712
net8711
net8710
net8709
net8708
net8707
net8706
net8705
net8704
net8703
net8702
net8701
net8700
net8699
net8698
net8697
net8696
net8695
net8694
net8693
net8692
net8691
net8690
net8689
net8688
net8687
net8686
net8685
net8684
net8683
net8682
net8681
net8680
net8679
net8678
net8677
net8676
net8675
net8674
net8673
net8672
net8671
net8670
net8669
net8668
net8667
net8666
net8665
net8664
net8663
net8662
net8661
net8660
net8659
net8658
net8657
net8656
net8655
net8654
net8653
net8652
net8651
net8650
net8649
net8648
net8647
net8646
net8645
net8644
net8643
net8642
net8641
net8640
net8639
net8638
net8637
net8636
net8635
net8633
net8632
net8631
net8630
net8629
net8627
net8626
net8625
net8624
net8623
net8622
net8621
net8620
net8619
net8618
net8617
net8616
net8615
net8614
net8613
net8612
net8611
net8610
net8609
net8608
net8607
net8606
net8605
net8604
net8603
net8602
net8601
net8600
net8599
net8598
net8597
net8596
net8595
net8594
net8593
net8592
net8591
net8590
net8589
net8588
net8587
net8586
net8585
net8584
net8583
net8582
net8581
net8580
net8579
net8578
net8577
net8576
net8575
net8574
net8573
net8572
net8571
net8570
net8569
net8568
net8567
net8566
net8565
net8564
net8563
net8562
net8561
net8560
net8559
net8558
net8557
net8556
net8555
net8554
net8553
net8552
net8551
net8550
net8549
net8548
net8547
net8546
net8545
net8544
net8543
net8542
net8541
net8540
net8539
net8538
net8537
net8536
net8535
net8534
net8533
net8532
net8531
net8530
net8529
net8528
net8527
net8526
net8525
net8524
net8523
net8522
net8521
net8520
net8519
net8518
net8517
net8516
net8515
net8514
net8513
net8512
net8511
net8510
net8509
net8508
net8507
net8506
net8505
net8504
net8503
net8502
net8501
net8500
net8499
net8498
net8497
net8496
net8495
net8494
net8493
net8492
net8491
net8490
net8489
net8488
net8487
net8486
net8485
net8484
net8483
net8482
net8481
net8480
net8479
net8478
net8477
net8476
net8475
net8474
net8473
net8472
net8471
net8470
net8469
net8468
net8467
net8466
net8465
net8464
net8463
net8462
net8461
net8460
net8459
net8458
net8457
net8456
net8455
net8454
net8453
net8452
net8451
net8450
net8449
net8448
net8447
net8446
net8445
net8444
net8443
net8442
net8441
net8440
net8439
net8438
net8437
net8436
net8435
net8434
net8433
net8432
net8431
net8430
net8429
net8427
net8426
net8425
net8424
net8423
net8422
net8421
net8420
net8419
net8418
net8417
net8416
net8415
net8414
net8413
net8412
net8411
net8410
net8409
net8408
net8407
net8406
net8405
net8404
net8403
net8402
net8401
net8400
net8399
net8398
net8397
net8396
net8395
net8394
net8393
net8392
net8391
net8390
net8389
net8388
net8387
net8386
net8385
net8384
net8383
net8382
net8381
net8380
net8379
net8378
net8377
net8376
net8375
net8374
net8373
net8372
net8371
net8370
net8369
net8368
net8367
net8366
net8365
net8364
net8363
net8362
net8361
net8360
net8359
net8358
net8357
net8356
net8355
net8354
net8353
net8352
net8351
net8350
net8349
net8348
net8347
net8346
net8345
net8344
net8343
net8342
net8341
net8340
net8339
net8338
net8337
net8336
net8335
net8334
net8333
net8332
net8331
net8330
net8329
net8328
net8327
net8326
net8325
net8324
net8323
net8322
net8321
net8320
net8319
net8318
net8317
net8316
net8315
net8314
net8313
net8312
net8311
net8310
net8309
net8308
net8307
net8306
net8305
net8304
net8303
net8302
net8301
net8300
net8299
net8298
net8297
net8296
net8295
net8294
net8293
net8292
net8291
net8290
net8289
net8288
net8287
net8286
net8285
net8284
net8283
net8282
net8281
net8280
net8279
net8278
net8277
net8276
net8275
net8274
net8273
net8272
net8271
net8270
net8269
net8268
net8267
net8266
net8265
net8264
net8263
net8262
net8261
net8260
net8259
net8258
net8257
net8256
net8255
net8254
net8253
net8252
net8251
net8250
net8249
net8248
net8247
net8246
net8245
net8244
net8243
net8242
net8241
net8240
net8239
net8238
net8237
net8236
net8235
net8234
net8233
net8232
net8231
net8230
net8229
net8228
net8227
net8226
net8225
net8224
net8223
net8222
net8221
net8220
net8219
net8218
net8217
net8216
net8215
net8214
net8213
net8212
net8211
net8210
net8209
net8208
net8207
net8206
net8205
net8204
net8203
net8202
net8201
net8200
net8199
net8198
net8197
net8196
net8195
net8194
net8193
net8192
net8191
net8190
net8189
net8188
net8187
net8186
net8185
net8184
net8183
net8182
net8181
net8180
net8179
net8178
net8177
net8176
net8175
net8174
net8173
net8172
net8171
net8170
net8169
net8168
net8167
net8166
net8165
net8164
net8163
net8162
net8161
net8160
net8159
net8158
net8157
net8156
net8155
net8154
net8153
net8152
net8151
net8150
net8149
net8148
net8147
net8146
net8145
net8144
net8143
net8142
net8141
net8140
net8139
net8138
net8137
net8136
net8135
net8134
net8133
net8132
net8131
net8130
net8129
net8128
net8127
net8126
net8125
net8124
net8123
net8122
net8121
net8120
net8119
net8118
net8117
net8116
net8115
net8114
net8113
net8112
net8111
net8110
net8109
net8108
net8107
net8106
net8105
net8104
net8103
net8102
net8101
net8100
net8099
net8097
net8096
net8095
net8094
net8093
net8092
net8091
net8090
net8089
net8088
net8087
net8086
net8085
net8084
net8083
net8082
net8081
net8080
net8079
net8078
net8077
net8076
net8075
net8074
net8073
net8072
net8071
net8070
net8069
net8068
net8067
net8066
net8065
net8064
net8063
net8062
net8061
net8060
net8059
net8058
net8057
net8056
net8055
net8054
net8053
net8052
net8051
net8050
net8049
net8048
net8047
net8046
net8045
net8044
net8043
net8042
net8041
net8040
net8039
net8038
net8037
net8036
net8035
net8034
net8033
net8032
net8031
net8030
net8029
net8028
net8027
net8026
net8025
net8024
net8023
net8022
net8021
net8020
net8019
net8018
net8017
net8016
net8015
net8014
net8013
net8012
net8011
net8010
net8009
net8008
net8007
net8006
net8005
net8004
net8003
net8002
net8001
net8000
net7999
net7998
net7997
net7996
net7995
net7994
net7993
net7992
net7991
net7990
net7989
net7988
net7987
net7986
net7985
net7984
net7983
net7982
net7981
net7980
net7979
net7978
net7977
net7976
net7975
net7974
net7973
net7972
net7971
net7970
net7969
net7967
net7966
net7965
net7964
net7963
net7962
net7961
net7960
net7959
net7958
net7957
net7956
net7955
net7954
net7953
net7952
net7951
net7950
net7949
net7948
net7947
net7946
net7945
net7944
net7943
net7942
net7941
net7940
net7939
net7938
net7937
net7936
net7935
net7934
net7933
net7932
net7931
net7930
net7929
net7928
net7927
net7926
net7925
net7924
net7923
net7922
net7921
net7920
net7919
net7918
net7917
net7916
net7915
net7914
net7913
net7912
net7911
net7910
net7909
net7908
net7907
net7906
net7905
net7904
net7903
net7902
net7901
net7900
net7899
net7898
net7897
net7896
net7895
net7894
net7893
net7892
net7891
net7890
net7889
net7888
net7887
net7886
net7885
net7884
net7883
net7882
net7881
net7880
net7879
net7878
net7877
net7876
net7875
net7874
net7873
net7872
net7871
net7870
net7869
net7868
net7867
net7866
net7865
net7864
net7863
net7862
net7861
net7860
net7859
net7858
net7857
net7856
net7855
net7854
net7853
net7852
net7851
net7850
net7849
net7848
net7847
net7846
net7845
net7844
net7843
net7842
net7841
net7840
net7839
net7838
net7837
net7836
net7835
net7834
net7833
net7832
net7831
net7830
net7829
net7828
net7827
net7826
net7825
net7824
net7823
net7822
net7821
net7820
net7819
net7818
net7817
net7816
net7815
net7814
net7813
net7812
net7811
net7810
net7809
net7808
net7807
net7806
net7805
net7804
net7803
net7802
net7801
net7800
net7799
net7798
net7797
net7796
net7795
net7794
net7793
net7792
net7791
net7790
net7789
net7788
net7787
net7786
net7785
net7784
net7783
net7782
net7781
net7780
net7779
net7778
net7777
net7776
net7775
net7774
net7773
net7771
net7770
net7769
net7768
net7767
net7766
net7765
net7764
net7763
net7762
net7761
net7760
net7759
net7758
net7757
net7756
net7755
net7754
net7753
net7752
net7751
net7750
net7749
net7748
net7747
net7746
net7745
net7744
net7743
net7742
net7741
net7740
net7739
net7738
net7737
net7736
net7735
net7734
net7733
net7732
net7731
net7730
net7729
net7728
net7727
net7726
net7725
net7724
net7723
net7722
net7721
net7720
net7719
net7718
net7717
net7716
net7715
net7714
net7713
net7712
net7711
net7710
net7709
net7708
net7707
net7706
net7705
net7704
net7703
net7702
net7700
net7699
net7698
net7697
net7696
net7695
net7694
net7693
net7692
net7691
net7690
net7689
net7688
net7687
net7686
net7685
net7684
net7683
net7682
net7681
net7680
net7679
net7678
net7677
net7676
net7675
net7674
net7673
net7672
net7671
net7670
net7669
net7668
net7667
net7666
net7665
net7664
net7663
net7662
net7661
net7660
net7659
net7658
net7657
net7656
net7655
net7654
net7653
net7652
net7651
net7650
net7648
net7647
net7646
net7645
net7644
net7643
net7642
net7641
net7640
net7639
net7638
net7637
net7636
net7635
net7634
net7633
net7632
net7631
net7630
net7629
net7627
net7626
net7625
net7624
net7623
net7622
net7621
net7620
net7619
net7618
net7617
net7616
net7615
net7614
net7613
net7612
net7611
net7610
net7609
net7608
net7607
net7606
net7605
net7604
net7603
net7602
net7601
net7600
net7599
net7598
net7597
net7596
net7595
net7594
net7593
net7592
net7591
net7590
net7589
net7588
net7587
net7586
net7585
net7584
net7583
net7582
net7581
net7580
net7579
net7578
net7577
net7576
net7575
net7574
net7573
net7572
net7571
net7570
net7569
net7568
net7567
net7566
net7565
net7564
net7562
net7561
net7560
net7559
net7558
net7557
net7556
net7555
net7554
net7553
net7552
net7551
net7550
net7549
net7548
net7547
net7546
net7545
net7544
net7543
net7542
net7541
net7540
net7539
net7538
net7536
net7535
net7534
net7533
net7532
net7531
net7530
net7529
net7528
net7527
net7526
net7525
net7524
net7523
net7522
net7521
net7520
net7519
net7518
net7517
net7516
net7515
net7514
net7513
net7512
net7511
net7510
net7509
net7508
net7507
net7506
net7505
net7504
net7503
net7502
net7501
net7500
net7499
net7498
net7497
net7496
net7495
net7494
net7493
net7492
net7491
net7490
net7489
net7488
net7487
net7486
net7485
net7484
net7483
net7482
net7481
net7480
net7479
net7478
net7477
net7476
net7475
net7474
net7473
net7472
net7471
net7470
net7469
net7468
net7467
net7466
net7465
net7464
net7463
net7462
net7461
net7460
net7459
net7458
net7457
net7456
net7455
net7454
net7453
net7452
net7451
net7450
net7449
net7448
net7447
net7446
net7445
net7444
net7443
net7442
net7441
net7440
net7439
net7437
net7436
net7435
net7434
net7433
net7432
net7431
net7430
net7429
net7428
net7427
net7426
net7425
net7424
net7423
net7422
net7421
net7420
net7419
net7418
net7417
net7416
net7415
net7414
net7413
net7412
net7411
net7410
net7409
net7408
net7407
net7406
net7405
net7404
net7403
net7402
net7401
net7400
net7399
net7398
net7397
net7396
net7395
net7394
net7393
net7392
net7391
net7390
net7389
net7388
net7387
net7386
net7385
net7384
net7383
net7382
net7381
net7380
net7379
net7378
net7377
net7376
net7375
net7374
net7373
net7372
net7371
net7370
net7369
net7368
net7367
net7366
net7365
net7364
net7363
net7362
net7361
net7360
net7359
net7358
net7357
net7356
net7355
net7354
net7353
net7352
net7351
net7350
net7349
net7348
net7347
net7346
net7345
net7344
net7343
net7342
net7341
net7340
net7339
net7338
net7337
net7336
net7335
net7334
net7333
net7332
net7331
net7330
net7329
net7328
net7327
net7326
net7325
net7324
net7322
net7321
net7320
net7319
net7318
net7317
net7316
net7315
net7314
net7313
net7312
net7310
net7309
net7308
net7307
net7306
net7305
net7304
net7303
net7302
net7301
net7300
net7299
net7298
net7297
net7296
net7295
net7294
net7293
net7292
net7291
net7290
net7289
net7288
net7287
net7286
net7285
net7284
net7283
net7282
net7281
net7280
net7279
net7278
net7277
net7276
net7275
net7274
net7273
net7272
net7271
net7270
net7269
net7268
net7267
net7266
net7265
net7264
net7263
net7262
net7261
net7260
net7259
net7258
net7257
net7256
net7255
net7254
net7253
net7252
net7251
net7250
net7249
net7248
net7247
net7246
net7245
net7244
net7243
net7242
net7241
net7240
net7239
net7238
net7237
net7236
net7235
net7234
net7233
net7232
net7231
net7230
net7229
net7228
net7227
net7226
net7225
net7224
net7223
net7222
net7221
net7220
net7219
net7218
net7217
net7216
net7215
net7214
net7213
net7212
net7211
net7210
net7209
net7208
net7207
net7206
net7205
net7204
net7203
net7202
net7201
net7200
net7199
net7198
net7197
net7196
net7195
net7194
net7193
net7192
net7191
net7190
net7189
net7188
net7187
net7186
net7185
net7184
net7183
net7182
net7181
net7180
net7179
net7178
net7177
net7176
net7175
net7174
net7173
net7172
net7171
net7170
net7169
net7168
net7167
net7166
net7165
net7164
net7163
net7162
net7161
net7160
net7159
net7158
net7157
net7156
net7155
net7154
net7153
net7152
net7151
net7150
net7149
net7148
net7147
net7146
net7145
net7144
net7143
net7142
net7141
net7140
net7139
net7138
net7137
net7136
net7135
net7134
net7133
net7132
net7131
net7130
net7129
net7128
net7127
net7126
net7125
net7124
net7123
net7122
net7121
net7120
net7119
net7118
net7117
net7116
net7115
net7114
net7113
net7112
net7111
net7110
net7109
net7108
net7107
net7106
net7105
net7104
net7103
net7102
net7101
net7100
net7099
net7098
net7097
net7096
net7095
net7094
net7093
net7092
net7091
net7090
net7089
net7088
net7087
net7086
net7085
net7084
net7083
net7082
net7081
net7080
net7079
net7078
net7077
net7076
net7075
net7074
net7073
net7072
net7071
net7070
net7069
net7068
net7067
net7066
net7065
net7064
net7063
net7062
net7061
net7060
net7059
net7058
net7057
net7056
net7055
net7054
net7053
net7052
net7051
net7050
net7049
net7048
net7047
net7046
net7045
net7044
net7043
net7042
net7041
net7040
net7039
net7038
net7037
net7036
net7035
net7034
net7033
net7032
net7031
net7030
net7029
net7028
net7027
net7025
net7024
net7023
net7022
net7021
net7020
net7019
net7018
net7017
net7016
net7015
net7014
net7013
net7012
net7011
net7010
net7009
net7008
net7007
net7006
net7005
net7003
net7002
net7001
net7000
net6999
net6998
net6997
net6996
net6995
net6994
net6993
net6992
net6991
net6990
net6989
net6988
net6987
net6986
net6985
net6984
net6983
net6982
net6981
net6980
net6979
net6978
net6977
net6976
net6975
net6974
net6973
net6972
net6971
net6970
net6969
net6968
net6967
net6966
net6965
net6964
net6963
net6962
net6961
net6960
net6959
net6958
net6957
net6956
net6955
net6954
net6953
net6952
net6951
net6950
net6949
net6948
net6947
net6946
net6945
net6944
net6943
net6942
net6941
net6940
net6939
net6938
net6937
net6936
net6935
net6934
net6933
net6932
net6931
net6930
net6929
net6928
net6927
net6926
net6925
net6924
net6923
net6922
net6921
net6920
net6919
net6918
net6917
net6916
net6915
net6914
net6913
net6912
net6911
net6910
net6909
net6908
net6907
net6906
net6905
net6904
net6903
net6902
net6901
net6900
net6899
net6898
net6897
net6896
net6895
net6894
net6893
net6892
net6891
net6890
net6889
net6888
net6887
net6886
net6885
net6884
net6883
net6882
net6881
net6880
net6879
net6878
net6877
net6876
net6875
net6874
net6873
net6872
net6871
net6870
net6869
net6868
net6867
net6866
net6865
net6864
net6863
net6862
net6861
net6860
net6859
net6858
net6857
net6855
net6854
net6853
net6852
net6851
net6850
net6849
net6848
net6847
net6846
net6845
net6844
net6843
net6842
net6841
net6840
net6839
net6838
net6837
net6836
net6835
net6834
net6833
net6832
net6831
net6830
net6829
net6828
net6827
net6826
net6825
net6824
net6823
net6822
net6820
net6819
net6818
net6817
net6816
net6815
net6814
net6813
net6812
net6811
net6810
net6809
net6808
net6807
net6806
net6805
net6804
net6803
net6802
net6801
net6800
net6799
net6798
net6797
net6795
net6794
net6793
net6792
net6791
net6790
net6789
net6788
net6787
net6786
net6785
net6784
net6783
net6782
net6781
net6780
net6779
net6778
net6777
net6776
net6775
net6774
net6773
net6772
net6771
net6770
net6769
net6768
net6767
net6766
net6765
net6764
net6763
net6762
net6761
net6760
net6759
net6758
net6757
net6756
net6755
net6754
net6753
net6752
net6751
net6750
net6749
net6748
net6747
net6746
net6745
net6744
net6743
net6742
net6741
net6740
net6739
net6738
net6737
net6736
net6735
net6734
net6733
net6732
net6731
net6730
net6729
net6728
net6727
net6726
net6725
net6724
net6723
net6722
net6721
net6720
net6719
net6718
net6717
net6716
net6715
net6714
net6713
net6712
net6711
net6710
net6709
net6708
net6707
net6706
net6705
net6704
net6703
net6702
net6701
net6700
net6699
net6698
net6697
net6696
net6695
net6694
net6693
net6692
net6691
net6690
net6689
net6688
net6687
net6686
net6685
net6684
net6683
net6682
net6681
net6680
net6679
net6678
net6677
net6676
net6675
net6674
net6673
net6672
net6671
net6670
net6669
net6668
net6667
net6666
net6665
net6664
net6663
net6662
net6661
net6660
net6659
net6658
net6656
net6655
net6654
net6653
net6652
net6651
net6650
net6649
net6648
net6647
net6646
net6645
net6644
net6643
net6642
net6641
net6640
net6639
net6638
net6637
net6636
net6635
net6634
net6633
net6632
net6631
net6630
net6629
net6628
net6627
net6626
net6625
net6624
net6623
net6622
net6621
net6620
net6619
net6618
net6617
net6616
net6615
net6614
net6613
net6612
net6611
net6610
net6609
net6608
net6607
net6606
net6605
net6604
net6603
net6602
net6601
net6600
net6599
net6598
net6597
net6596
net6595
net6594
net6593
net6592
net6591
net6590
net6589
net6588
net6587
net6586
net6585
net6584
net6583
net6582
net6581
net6580
net6579
net6578
net6577
net6576
net6575
net6574
net6573
net6572
net6571
net6570
net6569
net6568
net6567
net6566
net6565
net6564
net6563
net6562
net6561
net6560
net6559
net6558
net6557
net6556
net6555
net6554
net6553
net6552
net6551
net6549
net6548
net6547
net6546
net6545
net6544
net6543
net6542
net6541
net6540
net6539
net6538
net6537
net6536
net6535
net6534
net6533
net6532
net6531
net6530
net6529
net6528
net6527
net6526
net6525
net6524
net6523
net6522
net6521
net6520
net6519
net6518
net6517
net6516
net6515
net6514
net6513
net6512
net6511
net6510
net6509
net6508
net6507
net6506
net6505
net6504
net6503
net6502
net6501
net6500
net6499
net6498
net6497
net6496
net6495
net6494
net6493
net6492
net6491
net6490
net6489
net6488
net6487
net6486
net6485
net6484
net6483
net6482
net6481
net6480
net6479
net6478
net6477
net6476
net6475
net6474
net6473
net6472
net6471
net6470
net6469
net6468
net6467
net6466
net6465
net6464
net6463
net6462
net6461
net6460
net6459
net6458
net6457
net6456
net6455
net6454
net6453
net6452
net6451
net6450
net6449
net6448
net6447
net6446
net6445
net6444
net6443
net6442
net6441
net6440
net6439
net6438
net6437
net6436
net6435
net6434
net6433
net6431
net6430
net6429
net6428
net6427
net6426
net6425
net6424
net6423
net6422
net6421
net6420
net6419
net6418
net6417
net6416
net6415
net6414
net6413
net6412
net6411
net6410
net6409
net6408
net6407
net6406
net6405
net6404
net6403
net6402
net6401
net6400
net6399
net6398
net6397
net6396
net6395
net6394
net6393
net6392
net6391
net6390
net6389
net6388
net6387
net6386
net6385
net6384
net6383
net6382
net6381
net6380
net6379
net6378
net6377
net6376
net6375
net6374
net6373
net6372
net6371
net6370
net6369
net6368
net6367
net6366
net6365
net6364
net6363
net6362
net6361
net6360
net6359
net6358
net6357
net6356
net6355
net6354
net6353
net6352
net6351
net6350
net6349
net6348
net6347
net6346
net6345
net6344
net6343
net6342
net6341
net6340
net6339
net6338
net6337
net6336
net6335
net6334
net6333
net6332
net6331
net6330
net6329
net6328
net6327
net6326
net6325
net6324
net6323
net6322
net6321
net6320
net6319
net6318
net6317
net6316
net6315
net6314
net6313
net6312
net6311
net6310
net6309
net6308
net6307
net6306
net6305
net6304
net6303
net6302
net6301
net6300
net6299
net6298
net6297
net6296
net6295
net6294
net6293
net6292
net6291
net6290
net6289
net6288
net6287
net6286
net6285
net6284
net6283
net6282
net6281
net6280
net6279
net6278
net6277
net6276
net6275
net6274
net6273
net6272
net6271
net6270
net6269
net6268
net6267
net6266
net6265
net6264
net6263
net6262
net6261
net6260
net6259
net6258
net6257
net6256
net6255
net6254
net6253
net6252
net6251
net6250
net6249
net6248
net6247
net6246
net6245
net6244
net6243
net6242
net6241
net6240
net6239
net6238
net6237
net6236
net6235
net6234
net6233
net6232
net6231
net6230
net6229
net6228
net6227
net6226
net6225
net6224
net6223
net6222
net6221
net6220
net6219
net6218
net6217
net6216
net6215
net6214
net6213
net6212
net6211
net6210
net6209
net6208
net6207
net6206
net6205
net6204
net6203
net6202
net6201
net6200
net6199
net6198
net6197
net6196
net6195
net6194
net6193
net6192
net6191
net6190
net6189
net6188
net6187
net6186
net6185
net6184
net6183
net6182
net6181
net6180
net6179
net6178
net6177
net6175
net6174
net6173
net6172
net6171
net6170
net6169
net6168
net6167
net6166
net6165
net6164
net6163
net6162
net6161
net6160
net6159
net6158
net6157
net6156
net6155
net6154
net6153
net6152
net6151
net6150
net6149
net6148
net6147
net6146
net6145
net6144
net6143
net6142
net6141
net6140
net6139
net6138
net6137
net6136
net6135
net6134
net6132
net6131
net6130
net6129
net6128
net6127
net6126
net6125
net6124
net6123
net6122
net6121
net6120
net6119
net6118
net6117
net6116
net6115
net6114
net6113
net6112
net6111
net6110
net6109
net6108
net6106
net6105
net6104
net6103
net6102
net6101
net6100
net6099
net6098
net6097
net6096
net6095
net6094
net6093
net6092
net6091
net6090
net6089
net6088
net6087
net6086
net6085
net6084
net6083
net6082
net6081
net6080
net6079
net6078
net6077
net6076
net6075
net6074
net6073
net6072
net6071
net6070
net6069
net6068
net6067
net6066
net6065
net6064
net6063
net6062
net6061
net6060
net6059
net6058
net6057
net6056
net6055
net6054
net6053
net6052
net6051
net6050
net6049
net6048
net6047
net6046
net6045
net6044
net6043
net6042
net6041
net6040
net6039
net6038
net6037
net6036
net6035
net6034
net6033
net6032
net6031
net6030
net6029
net6028
net6027
net6026
net6025
net6024
net6023
net6022
net6021
net6020
net6019
net6018
net6017
net6016
net6015
net6014
net6013
net6012
net6011
net6010
net6009
net6008
net6007
net6006
net6005
net6004
net6003
net6002
net6001
net6000
net5999
net5998
net5997
net5996
net5995
net5994
net5993
net5992
net5991
net5990
net5989
net5988
net5987
net5986
net5985
net5984
net5983
net5982
net5981
net5980
net5979
net5978
net5977
net5976
net5975
net5974
net5973
net5972
net5971
net5970
net5969
net5968
net5967
net5966
net5965
net5964
net5963
net5962
net5961
net5960
net5959
net5958
net5957
net5956
net5955
net5954
net5953
net5952
net5951
net5950
net5949
net5948
net5947
net5946
net5945
net5944
net5943
net5942
net5941
net5940
net5939
net5938
net5937
net5936
net5935
net5934
net5933
net5932
net5931
net5930
net5929
net5928
net5927
net5926
net5925
net5924
net5923
net5922
net5921
net5920
net5919
net5918
net5917
net5916
net5915
net5914
net5913
net5912
net5911
net5910
net5909
net5908
net5907
net5906
net5905
net5904
net5903
net5902
net5901
net5900
net5899
net5898
net5897
net5896
net5895
net5894
net5893
net5892
net5891
net5890
net5889
net5888
net5887
net5886
net5885
net5884
net5883
net5882
net5881
net5880
net5879
net5878
net5877
net5876
net5875
net5874
net5873
net5872
net5871
net5870
net5869
net5868
net5867
net5866
net5865
net5864
net5863
net5862
net5861
net5860
net5859
net5858
net5857
net5856
net5855
net5854
net5853
net5852
net5851
net5850
net5849
net5848
net5847
net5846
net5845
net5844
net5843
net5842
net5841
net5840
net5839
net5838
net5837
net5836
net5835
net5834
net5833
net5832
net5831
net5830
net5829
net5828
net5827
net5826
net5825
net5824
net5823
net5822
net5821
net5820
net5819
net5818
net5817
net5816
net5815
net5814
net5813
net5812
net5811
net5810
net5809
net5808
net5807
net5806
net5805
net5804
net5803
net5802
net5801
net5800
net5799
net5798
net5797
net5796
net5795
net5794
net5793
net5792
net5791
net5790
net5789
net5787
net5786
net5785
net5784
net5783
net5782
net5781
net5780
net5779
net5778
net5777
net5776
net5775
net5774
net5773
net5772
net5771
net5770
net5769
net5768
net5767
net5766
net5765
net5764
net5763
net5762
net5761
net5760
net5759
net5758
net5757
net5756
net5755
net5754
net5753
net5752
net5751
net5750
net5749
net5748
net5747
net5746
net5745
net5744
net5743
net5742
net5741
net5740
net5739
net5738
net5737
net5736
net5735
net5734
net5733
net5732
net5731
net5730
net5729
net5728
net5727
net5726
net5725
net5724
net5723
net5722
net5721
net5720
net5718
net5717
net5716
net5715
net5714
net5713
net5712
net5711
net5710
net5709
net5708
net5707
net5706
net5705
net5704
net5703
net5702
net5701
net5700
net5699
net5698
net5697
net5696
net5695
net5694
net5693
net5692
net5691
net5690
net5689
net5688
net5687
net5686
net5685
net5684
net5683
net5682
net5681
net5680
net5679
net5678
net5677
net5676
net5675
net5674
net5673
net5672
net5671
net5670
net5669
net5668
net5667
net5666
net5665
net5664
net5663
net5662
net5661
net5660
net5659
net5658
net5657
net5656
net5655
net5654
net5653
net5652
net5651
net5650
net5649
net5648
net5647
net5646
net5645
net5644
net5643
net5642
net5641
net5640
net5639
net5638
net5637
net5636
net5635
net5634
net5633
net5632
net5631
net5630
net5629
net5628
net5627
net5626
net5625
net5624
net5623
net5622
net5621
net5620
net5619
net5618
net5617
net5616
net5615
net5614
net5613
net5612
net5611
net5610
net5609
net5608
net5607
net5606
net5605
net5604
net5603
net5602
net5601
net5600
net5599
net5598
net5597
net5596
net5595
net5594
net5593
net5592
net5591
net5590
net5589
net5588
net5587
net5586
net5585
net5584
net5583
net5582
net5581
net5580
net5579
net5578
net5577
net5576
net5575
net5574
net5573
net5572
net5571
net5570
net5569
net5568
net5567
net5566
net5565
net5564
net5563
net5562
net5561
net5560
net5559
net5558
net5557
net5556
net5555
net5554
net5553
net5552
net5551
net5550
net5549
net5548
net5547
net5546
net5545
net5544
net5543
net5542
net5541
net5540
net5539
net5538
net5537
net5536
net5535
net5534
net5533
net5531
net5530
net5529
net5528
net5527
net5526
net5525
net5524
net5523
net5522
net5521
net5520
net5519
net5518
net5517
net5516
net5515
net5514
net5513
net5512
net5511
net5510
net5509
net5508
net5507
net5506
net5505
net5504
net5503
net5502
net5501
net5500
net5499
net5498
net5497
net5496
net5495
net5494
net5493
net5492
net5491
net5490
net5489
net5488
net5487
net5486
net5485
net5484
net5483
net5482
net5481
net5480
net5479
net5478
net5477
net5476
net5475
net5474
net5473
net5472
net5471
net5470
net5469
net5468
net5467
net5466
net5465
net5464
net5463
net5462
net5461
net5460
net5459
net5458
net5457
net5456
net5455
net5454
net5453
net5452
net5451
net5450
net5449
net5448
net5447
net5446
net5445
net5444
net5443
net5442
net5441
net5440
net5439
net5438
net5437
net5436
net5435
net5434
net5433
net5432
net5431
net5430
net5429
net5428
net5427
net5426
net5425
net5424
net5423
net5422
net5421
net5420
net5419
net5418
net5417
net5416
net5415
net5414
net5413
net5412
net5411
net5410
net5409
net5408
net5407
net5406
net5405
net5404
net5403
net5402
net5401
net5400
net5399
net5398
net5397
net5396
net5395
net5394
net5393
net5392
net5391
net5390
net5389
net5388
net5387
net5386
net5385
net5384
net5383
net5381
net5380
net5379
net5378
net5377
net5376
net5375
net5374
net5373
net5372
net5371
net5370
net5369
net5368
net5367
net5366
net5365
net5364
net5363
net5362
net5361
net5360
net5359
net5358
net5357
net5356
net5355
net5354
net5353
net5352
net5351
net5350
net5349
net5348
net5347
net5346
net5345
net5344
net5343
net5342
net5341
net5340
net5339
net5338
net5337
net5336
net5335
net5334
net5333
net5332
net5331
net5330
net5329
net5328
net5327
net5326
net5325
net5324
net5323
net5322
net5321
net5320
net5319
net5318
net5317
net5316
net5315
net5314
net5313
net5312
net5311
net5310
net5309
net5308
net5307
net5306
net5305
net5304
net5303
net5302
net5301
net5300
net5299
net5298
net5297
net5296
net5295
net5294
net5293
net5292
net5291
net5290
net5289
net5288
net5287
net5286
net5285
net5284
net5283
net5282
net5281
net5280
net5279
net5278
net5277
net5276
net5275
net5274
net5273
net5272
net5271
net5270
net5269
net5268
net5267
net5266
net5265
net5264
net5263
net5262
net5261
net5260
net5259
net5258
net5257
net5256
net5255
net5254
net5253
net5252
net5251
net5250
net5249
net5248
net5247
net5246
net5245
net5244
net5243
net5242
net5241
net5240
net5239
net5238
net5237
net5236
net5235
net5234
net5233
net5232
net5231
net5230
net5229
net5228
net5227
net5226
net5225
net5224
net5223
net5222
net5221
net5220
net5219
net5218
net5217
net5216
net5215
net5214
net5213
net5212
net5211
net5210
net5209
net5208
net5207
net5206
net5205
net5204
net5203
net5202
net5201
net5200
net5199
net5198
net5197
net5196
net5195
net5194
net5193
net5192
net5191
net5190
net5189
net5188
net5187
net5186
net5185
net5184
net5183
net5182
net5181
net5180
net5179
net5178
net5177
net5176
net5175
net5174
net5173
net5172
net5171
net5170
net5169
net5168
net5167
net5166
net5165
net5164
net5163
net5162
net5161
net5160
net5159
net5158
net5157
net5156
net5155
net5154
net5153
net5152
net5151
net5150
net5149
net5148
net5147
net5146
net5145
net5144
net5143
net5142
net5141
net5140
net5139
net5138
net5137
net5136
net5135
net5134
net5133
net5132
net5131
net5130
net5129
net5128
net5127
net5126
net5125
net5124
net5123
net5122
net5121
net5120
net5119
net5118
net5117
net5116
net5115
net5114
net5113
net5112
net5111
net5110
net5109
net5108
net5107
net5106
net5105
net5104
net5103
net5102
net5101
net5100
net5099
net5098
net5097
net5096
net5095
net5094
net5093
net5092
net5091
net5090
net5089
net5088
net5087
net5086
net5085
net5084
net5083
net5082
net5081
net5080
net5079
net5078
net5077
net5076
net5075
net5073
net5072
net5071
net5070
net5069
net5068
net5067
net5066
net5065
net5064
net5063
net5062
net5061
net5060
net5059
net5058
net5057
net5056
net5055
net5054
net5053
net5052
net5051
net5050
net5049
net5048
net5047
net5046
net5045
net5044
net5043
net5042
net5041
net5040
net5039
net5038
net5037
net5036
net5035
net5034
net5033
net5032
net5031
net5030
net5029
net5028
net5027
net5026
net5025
net5024
net5023
net5022
net5020
net5019
net5018
net5017
net5016
net5015
net5014
net5013
net5012
net5011
net5010
net5009
net5008
net5007
net5006
net5005
net5004
net5003
net5002
net5001
net5000
net4999
net4998
net4997
net4996
net4995
net4994
net4993
net4992
net4991
net4990
net4989
net4988
net4987
net4986
net4985
net4984
net4983
net4982
net4981
net4980
net4979
net4978
net4977
net4976
net4975
net4974
net4973
net4972
net4971
net4970
net4969
net4968
net4967
net4966
net4965
net4964
net4963
net4962
net4961
net4960
net4959
net4958
net4957
net4956
net4955
net4954
net4953
net4952
net4951
net4950
net4949
net4948
net4947
net4946
net4945
net4944
net4943
net4942
net4941
net4940
net4939
net4938
net4937
net4936
net4935
net4934
net4933
net4932
net4931
net4930
net4929
net4928
net4927
net4926
net4925
net4924
net4923
net4922
net4921
net4920
net4919
net4918
net4917
net4916
net4915
net4914
net4913
net4912
net4911
net4910
net4909
net4908
net4907
net4906
net4905
net4904
net4903
net4902
net4901
net4900
net4899
net4898
net4897
net4896
net4895
net4894
net4893
net4892
net4891
net4890
net4889
net4888
net4887
net4886
net4885
net4884
net4883
net4882
net4881
net4880
net4879
net4878
net4877
net4876
net4875
net4874
net4873
net4872
net4871
net4870
net4869
net4868
net4867
net4866
net4865
net4864
net4863
net4862
net4861
net4860
net4859
net4858
net4857
net4856
net4855
net4854
net4853
net4852
net4851
net4850
net4849
net4848
net4847
net4846
net4845
net4844
net4843
net4842
net4841
net4840
net4839
net4838
net4837
net4836
net4835
net4834
net4833
net4832
net4831
net4830
net4829
net4828
net4827
net4826
net4825
net4824
net4823
net4822
net4821
net4820
net4819
net4818
net4817
net4816
net4815
net4814
net4813
net4812
net4811
net4810
net4809
net4808
net4807
net4806
net4805
net4804
net4803
net4802
net4801
net4800
net4799
net4798
net4797
net4796
net4794
net4793
net4792
net4791
net4790
net4789
net4788
net4787
net4786
net4785
net4784
net4783
net4782
net4781
net4780
net4779
net4778
net4777
net4776
net4775
net4774
net4773
net4772
net4771
net4770
net4769
net4768
net4767
net4766
net4765
net4764
net4763
net4762
net4761
net4760
net4759
net4758
net4757
net4756
net4755
net4754
net4753
net4752
net4751
net4750
net4749
net4748
net4747
net4746
net4745
net4744
net4743
net4742
net4741
net4740
net4739
net4738
net4737
net4736
net4735
net4734
net4733
net4732
net4731
net4730
net4729
net4728
net4727
net4726
net4725
net4724
net4723
net4722
net4721
net4720
net4719
net4718
net4717
net4716
net4715
net4714
net4713
net4712
net4711
net4710
net4709
net4708
net4707
net4706
net4705
net4704
net4703
net4702
net4701
net4700
net4699
net4698
net4697
net4696
net4695
net4694
net4693
net4692
net4691
net4690
net4689
net4688
net4687
net4686
net4685
net4684
net4682
net4681
net4680
net4679
net4678
net4677
net4676
net4675
net4674
net4673
net4672
net4671
net4670
net4669
net4668
net4667
net4666
net4665
net4664
net4663
net4662
net4661
net4660
net4659
net4658
net4657
net4656
net4655
net4654
net4653
net4652
net4651
net4650
net4649
net4648
net4647
net4646
net4645
net4644
net4643
net4642
net4641
net4640
net4639
net4638
net4637
net4636
net4635
net4634
net4633
net4632
net4630
net4629
net4628
net4627
net4626
net4625
net4624
net4623
net4622
net4621
net4620
net4619
net4618
net4617
net4616
net4615
net4614
net4613
net4612
net4611
net4610
net4609
net4608
net4607
net4606
net4605
net4604
net4603
net4602
net4601
net4600
net4599
net4598
net4597
net4596
net4595
net4594
net4593
net4592
net4591
net4590
net4589
net4588
net4587
net4586
net4585
net4584
net4583
net4582
net4581
net4580
net4579
net4578
net4577
net4576
net4575
net4574
net4573
net4572
net4571
net4570
net4569
net4568
net4567
net4566
net4565
net4564
net4563
net4562
net4561
net4560
net4559
net4558
net4557
net4556
net4555
net4554
net4553
net4552
net4551
net4550
net4549
net4548
net4547
net4546
net4545
net4544
net4543
net4542
net4541
net4540
net4539
net4538
net4537
net4536
net4535
net4534
net4533
net4532
net4531
net4530
net4529
net4528
net4527
net4526
net4525
net4524
net4523
net4522
net4521
net4520
net4519
net4518
net4517
net4516
net4515
net4514
net4513
net4512
net4511
net4510
net4509
net4508
net4507
net4506
net4505
net4504
net4503
net4501
net4500
net4499
net4498
net4497
net4496
net4495
net4494
net4493
net4492
net4491
net4490
net4489
net4488
net4487
net4486
net4485
net4484
net4483
net4482
net4481
net4480
net4479
net4478
net4477
net4476
net4475
net4474
net4473
net4472
net4471
net4470
net4469
net4468
net4467
net4466
net4465
net4464
net4463
net4462
net4461
net4460
net4459
net4458
net4457
net4456
net4455
net4454
net4453
net4452
net4451
net4450
net4449
net4448
net4447
net4446
net4445
net4444
net4443
net4442
net4441
net4440
net4439
net4438
net4437
net4436
net4435
net4434
net4433
net4432
net4431
net4430
net4429
net4428
net4427
net4426
net4425
net4424
net4423
net4422
net4421
net4420
net4419
net4418
net4417
net4416
net4415
net4414
net4413
net4412
net4411
net4410
net4409
net4408
net4407
net4406
net4405
net4404
net4403
net4402
net4401
net4400
net4399
net4398
net4397
net4396
net4395
net4394
net4393
net4392
net4391
net4390
net4389
net4388
net4387
net4386
net4385
net4384
net4383
net4382
net4381
net4380
net4379
net4378
net4377
net4376
net4375
net4374
net4373
net4372
net4371
net4370
net4369
net4368
net4367
net4366
net4365
net4364
net4363
net4362
net4361
net4360
net4359
net4358
net4357
net4356
net4355
net4354
net4353
net4352
net4351
net4350
net4349
net4348
net4347
net4346
net4345
net4344
net4343
net4342
net4341
net4340
net4339
net4338
net4337
net4336
net4335
net4334
net4333
net4332
net4331
net4330
net4329
net4328
net4327
net4326
net4325
net4324
net4323
net4322
net4321
net4320
net4319
net4318
net4317
net4316
net4315
net4314
net4313
net4312
net4311
net4310
net4309
net4308
net4307
net4306
net4305
net4304
net4303
net4302
net4301
net4300
net4299
net4298
net4297
net4296
net4295
net4294
net4293
net4292
net4291
net4290
net4289
net4288
net4287
net4286
net4285
net4284
net4283
net4282
net4281
net4280
net4279
net4278
net4277
net4276
net4275
net4274
net4273
net4272
net4271
net4270
net4269
net4268
net4267
net4266
net4265
net4263
net4262
net4261
net4260
net4259
net4258
net4257
net4256
net4255
net4254
net4253
net4252
net4251
net4250
net4249
net4248
net4247
net4246
net4245
net4244
net4243
net4242
net4241
net4240
net4238
net4237
net4236
net4235
net4234
net4233
net4232
net4231
net4230
net4229
net4228
net4227
net4226
net4225
net4224
net4223
net4222
net4221
net4220
net4219
net4218
net4217
net4216
net4215
net4214
net4213
net4212
net4211
net4210
net4209
net4208
net4207
net4206
net4205
net4204
net4203
net4202
net4201
net4200
net4199
net4198
net4197
net4196
net4195
net4194
net4193
net4192
net4191
net4190
net4189
net4188
net4187
net4186
net4185
net4184
net4183
net4182
net4181
net4180
net4179
net4178
net4177
net4176
net4175
net4174
net4173
net4172
net4171
net4170
net4169
net4168
net4167
net4166
net4165
net4164
net4163
net4162
net4161
net4160
net4159
net4158
net4157
net4156
net4155
net4154
net4153
net4152
net4151
net4150
net4149
net4148
net4147
net4146
net4145
net4144
net4143
net4142
net4141
net4140
net4139
net4138
net4137
net4136
net4135
net4134
net4133
net4132
net4131
net4130
net4129
net4128
net4127
net4126
net4125
net4124
net4123
net4122
net4121
net4120
net4119
net4118
net4117
net4116
net4115
net4114
net4113
net4112
net4111
net4110
net4109
net4108
net4107
net4106
net4105
net4104
net4103
net4102
net4101
net4100
net4099
net4098
net4097
net4096
net4095
net4094
net4093
net4092
net4091
net4090
net4089
net4088
net4087
net4086
net4085
net4084
net4083
net4082
net4081
net4080
net4079
net4078
net4077
net4076
net4075
net4074
net4073
net4072
net4071
net4070
net4069
net4068
net4067
net4066
net4065
net4064
net4063
net4062
net4061
net4060
net4059
net4058
net4056
net4055
net4054
net4053
net4052
net4051
net4050
net4049
net4048
net4047
net4046
net4045
net4044
net4043
net4042
net4041
net4040
net4039
net4038
net4037
net4036
net4035
net4034
net4033
net4032
net4031
net4030
net4029
net4028
net4027
net4026
net4025
net4024
net4023
net4022
net4021
net4020
net4019
net4018
net4017
net4016
net4015
net4014
net4013
net4012
net4011
net4010
net4009
net4008
net4007
net4006
net4005
net4004
net4003
net4002
net4001
net4000
net3999
net3998
net3997
net3996
net3995
net3994
net3993
net3992
net3991
net3990
net3989
net3988
net3987
net3986
net3985
net3984
net3983
net3982
net3981
net3980
net3979
net3978
net3977
net3976
net3975
net3974
net3973
net3972
net3971
net3970
net3969
net3968
net3967
net3966
net3965
net3964
net3963
net3962
net3961
net3960
net3959
net3958
net3957
net3956
net3955
net3954
net3953
net3952
net3951
net3950
net3949
net3948
net3946
net3945
net3944
net3943
net3942
net3941
net3940
net3939
net3938
net3937
net3936
net3935
net3934
net3933
net3932
net3931
net3930
net3929
net3928
net3927
net3926
net3925
net3924
net3923
net3922
net3921
net3920
net3919
net3918
net3917
net3916
net3915
net3914
net3913
net3912
net3911
net3910
net3909
net3908
net3907
net3906
net3905
net3904
net3903
net3902
net3901
net3900
net3899
net3898
net3897
net3896
net3895
net3894
net3893
net3892
net3891
net3890
net3889
net3888
net3887
net3886
net3885
net3884
net3883
net3882
net3881
net3880
net3879
net3878
net3877
net3876
net3875
net3874
net3873
net3872
net3871
net3870
net3869
net3868
net3867
net3866
net3865
net3864
net3863
net3862
net3861
net3860
net3859
net3858
net3857
net3856
net3855
net3854
net3853
net3852
net3851
net3850
net3849
net3848
net3847
net3846
net3845
net3844
net3843
net3842
net3841
net3840
net3839
net3838
net3837
net3836
net3835
net3834
net3833
net3832
net3831
net3830
net3829
net3828
net3827
net3826
net3825
net3824
net3823
net3822
net3821
net3820
net3819
net3818
net3817
net3816
net3815
net3814
net3813
net3812
net3811
net3810
net3809
net3808
net3807
net3806
net3805
net3804
net3803
net3802
net3801
net3800
net3799
net3798
net3797
net3796
net3795
net3794
net3793
net3792
net3791
net3790
net3789
net3788
net3787
net3786
net3785
net3784
net3783
net3782
net3781
net3780
net3779
net3778
net3777
net3776
net3775
net3774
net3773
net3772
net3771
net3770
net3769
net3768
net3767
net3766
net3765
net3764
net3763
net3762
net3761
net3760
net3759
net3758
net3757
net3756
net3755
net3754
net3753
net3752
net3751
net3750
net3749
net3748
net3747
net3746
net3745
net3744
net3743
net3742
net3741
net3740
net3739
net3738
net3737
net3736
net3735
net3734
net3733
net3732
net3731
net3730
net3729
net3728
net3727
net3726
net3725
net3724
net3723
net3722
net3721
net3720
net3719
net3718
net3717
net3716
net3715
net3714
net3713
net3712
net3711
net3710
net3709
net3708
net3707
net3706
net3705
net3704
net3703
net3702
net3701
net3700
net3699
net3698
net3697
net3696
net3695
net3694
net3693
net3692
net3691
net3690
net3689
net3688
net3687
net3686
net3685
net3684
net3683
net3682
net3681
net3680
net3679
net3678
net3677
net3676
net3675
net3674
net3673
net3672
net3671
net3670
net3669
net3668
net3667
net3666
net3665
net3664
net3663
net3662
net3661
net3660
net3659
net3658
net3657
net3656
net3655
net3654
net3653
net3652
net3651
net3650
net3649
net3648
net3647
net3646
net3645
net3644
net3643
net3642
net3641
net3640
net3639
net3638
net3637
net3636
net3635
net3634
net3633
net3632
net3631
net3630
net3629
net3628
net3627
net3626
net3625
net3624
net3623
net3622
net3621
net3620
net3619
net3618
net3617
net3616
net3615
net3614
net3613
net3612
net3611
net3610
net3609
net3608
net3607
net3606
net3605
net3604
net3603
net3602
net3601
net3600
net3599
net3598
net3597
net3596
net3595
net3594
net3593
net3592
net3591
net3590
net3589
net3588
net3587
net3586
net3585
net3584
net3582
net3581
net3580
net3579
net3578
net3577
net3576
net3575
net3574
net3573
net3572
net3571
net3570
net3569
net3568
net3567
net3566
net3565
net3564
net3563
net3562
net3561
net3560
net3559
net3558
net3557
net3556
net3555
net3554
net3553
net3552
net3551
net3550
net3549
net3548
net3547
net3546
net3545
net3544
net3543
net3542
net3541
net3540
net3539
net3538
net3537
net3536
net3535
net3534
net3533
net3532
net3531
net3530
net3529
net3528
net3527
net3526
net3525
net3524
net3523
net3522
net3521
net3520
net3519
net3518
net3517
net3516
net3515
net3514
net3513
net3512
net3511
net3510
net3509
net3508
net3507
net3506
net3505
net3504
net3503
net3502
net3501
net3500
net3499
net3498
net3497
net3496
net3495
net3494
net3493
net3492
net3491
net3490
net3489
net3488
net3487
net3486
net3485
net3484
net3483
net3482
net3481
net3480
net3479
net3478
net3477
net3476
net3475
net3474
net3473
net3472
net3471
net3470
net3469
net3468
net3467
net3466
net3465
net3464
net3463
net3462
net3461
net3460
net3459
net3458
net3457
net3456
net3455
net3454
net3453
net3452
net3451
net3450
net3449
net3448
net3447
net3446
net3445
net3444
net3443
net3442
net3441
net3440
net3439
net3438
net3437
net3436
net3435
net3434
net3433
net3432
net3431
net3430
net3429
net3428
net3427
net3426
net3425
net3424
net3423
net3422
net3421
net3420
net3419
net3418
net3417
net3416
net3415
net3414
net3413
net3412
net3411
net3410
net3409
net3408
net3407
net3406
net3405
net3404
net3403
net3402
net3401
net3400
net3399
net3398
net3397
net3396
net3395
net3394
net3393
net3392
net3391
net3390
net3389
net3388
net3387
net3386
net3385
net3384
net3383
net3382
net3381
net3380
net3379
net3378
net3377
net3376
net3375
net3374
net3373
net3372
net3371
net3370
net3369
net3368
net3367
net3366
net3365
net3364
net3363
net3362
net3361
net3360
net3359
net3358
net3357
net3356
net3355
net3354
net3353
net3352
net3351
net3350
net3349
net3348
net3347
net3346
net3345
net3344
net3343
net3342
net3341
net3340
net3339
net3338
net3337
net3336
net3335
net3334
net3333
net3332
net3331
net3330
net3329
net3328
net3327
net3326
net3325
net3324
net3323
net3322
net3321
net3320
net3319
net3318
net3317
net3316
net3315
net3314
net3313
net3312
net3311
net3310
net3309
net3308
net3307
net3306
net3305
net3304
net3303
net3302
net3301
net3300
net3299
net3298
net3297
net3296
net3295
net3294
net3293
net3292
net3291
net3290
net3289
net3288
net3287
net3286
net3285
net3284
net3283
net3282
net3281
net3280
net3279
net3278
net3277
net3276
net3275
net3274
net3273
net3272
net3271
net3270
net3269
net3268
net3267
net3266
net3265
net3264
net3263
net3262
net3261
net3260
net3259
net3258
net3257
net3256
net3255
net3254
net3253
net3252
net3251
net3250
net3249
net3248
net3247
net3246
net3245
net3244
net3243
net3242
net3241
net3240
net3239
net3238
net3237
net3236
net3235
net3234
net3233
net3232
net3231
net3230
net3229
net3228
net3227
net3226
net3225
net3224
net3223
net3222
net3221
net3220
net3219
net3218
net3217
net3216
net3215
net3214
net3213
net3212
net3211
net3210
net3209
net3208
net3207
net3206
net3205
net3204
net3203
net3202
net3201
net3200
net3199
net3198
net3197
net3196
net3195
net3194
net3193
net3192
net3191
net3190
net3189
net3188
net3187
net3186
net3185
net3184
net3183
net3182
net3181
net3180
net3179
net3178
net3177
net3176
net3175
net3174
net3173
net3172
net3171
net3170
net3169
net3168
net3167
net3166
net3165
net3164
net3163
net3161
net3160
net3159
net3158
net3157
net3156
net3155
net3154
net3153
net3152
net3151
net3150
net3149
net3148
net3147
net3146
net3145
net3144
net3143
net3142
net3141
net3140
net3139
net3138
net3137
net3136
net3135
net3134
net3133
net3132
net3131
net3130
net3129
net3128
net3127
net3126
net3125
net3124
net3123
net3122
net3121
net3120
net3119
net3118
net3117
net3116
net3115
net3114
net3113
net3112
net3111
net3110
net3109
net3108
net3107
net3106
net3105
net3104
net3103
net3102
net3101
net3100
net3099
net3098
net3097
net3096
net3095
net3094
net3093
net3092
net3091
net3090
net3089
net3088
net3087
net3086
net3085
net3084
net3083
net3082
net3081
net3080
net3079
net3078
net3077
net3076
net3075
net3074
net3073
net3072
net3071
net3070
net3069
net3068
net3067
net3066
net3065
net3064
net3063
net3062
net3061
net3060
net3059
net3058
net3057
net3056
net3055
net3054
net3053
net3052
net3051
net3050
net3049
net3048
net3047
net3046
net3045
net3044
net3043
net3042
net3041
net3040
net3039
net3038
net3037
net3036
net3035
net3034
net3033
net3032
net3031
net3030
net3029
net3028
net3027
net3026
net3025
net3024
net3023
net3022
net3021
net3020
net3019
net3018
net3017
net3016
net3015
net3014
net3013
net3012
net3011
net3010
net3009
net3008
net3007
net3006
net3005
net3004
net3003
net3002
net3001
net3000
net2999
net2998
net2997
net2996
net2995
net2994
net2993
net2992
net2991
net2990
net2989
net2988
net2987
net2986
net2985
net2984
net2983
net2982
net2981
net2980
net2979
net2978
net2977
net2976
net2975
net2974
net2973
net2972
net2971
net2970
net2969
net2968
net2967
net2966
net2965
net2964
net2963
net2962
net2961
net2960
net2959
net2958
net2957
net2956
net2955
net2954
net2953
net2952
net2951
net2950
net2949
net2948
net2947
net2946
net2945
net2944
net2943
net2942
net2941
net2940
net2939
net2938
net2937
net2936
net2935
net2934
net2933
net2932
net2931
net2930
net2929
net2928
net2927
net2926
net2925
net2924
net2923
net2922
net2921
net2920
net2919
net2918
net2917
net2916
net2915
net2914
net2913
net2912
net2911
net2910
net2909
net2908
net2907
net2906
net2905
net2904
net2903
net2902
net2901
net2900
net2899
net2898
net2897
net2896
net2895
net2894
net2893
net2892
net2891
net2890
net2889
net2888
net2887
net2886
net2885
net2884
net2883
net2882
net2881
net2880
net2879
net2878
net2877
net2876
net2875
net2874
net2873
net2872
net2871
net2870
net2869
net2868
net2867
net2866
net2865
net2864
net2863
net2862
net2861
net2860
net2859
net2858
net2857
net2856
net2855
net2854
net2853
net2852
net2851
net2850
net2849
net2848
net2847
net2846
net2845
net2844
net2843
net2842
net2841
net2840
net2839
net2838
net2837
net2836
net2835
net2834
net2833
net2832
net2831
net2830
net2829
net2828
net2827
net2826
net2825
net2824
net2823
net2822
net2821
net2820
net2819
net2818
net2817
net2816
net2815
net2814
net2813
net2812
net2811
net2810
net2809
net2808
net2807
net2806
net2805
net2804
net2803
net2802
net2801
net2800
net2799
net2798
net2797
net2796
net2795
net2794
net2793
net2792
net2791
net2790
net2789
net2788
net2787
net2786
net2785
net2784
net2783
net2782
net2781
net2780
net2779
net2778
net2777
net2776
net2775
net2774
net2773
net2772
net2771
net2770
net2769
net2768
net2767
net2766
net2765
net2764
net2763
net2762
net2761
net2760
net2759
net2758
net2757
net2756
net2755
net2754
net2753
net2752
net2751
net2750
net2749
net2748
net2747
net2746
net2745
net2744
net2743
net2742
net2741
net2740
net2739
net2738
net2737
net2736
net2735
net2734
net2733
net2732
net2731
net2730
net2729
net2728
net2727
net2726
net2725
net2724
net2723
net2722
net2721
net2720
net2719
net2718
net2717
net2716
net2715
net2714
net2713
net2712
net2711
net2710
net2709
net2708
net2707
net2706
net2705
net2704
net2703
net2702
net2701
net2700
net2699
net2698
net2697
net2696
net2695
net2694
net2693
net2692
net2691
net2690
net2689
net2688
net2687
net2686
net2685
net2684
net2683
net2682
net2681
net2680
net2679
net2678
net2677
net2676
net2675
net2674
net2673
net2672
net2671
net2670
net2669
net2668
net2667
net2666
net2665
net2664
net2663
net2662
net2661
net2660
net2659
net2658
net2657
net2656
net2655
net2654
net2653
net2652
net2651
net2650
net2648
net2647
net2646
net2645
net2644
net2643
net2642
net2641
net2640
net2639
net2638
net2637
net2636
net2635
net2634
net2633
net2632
net2631
net2630
net2629
net2628
net2627
net2626
net2625
net2624
net2623
net2622
net2621
net2620
net2619
net2618
net2617
net2616
net2615
net2614
net2613
net2612
net2611
net2610
net2609
net2608
net2607
net2606
net2605
net2604
net2603
net2602
net2601
net2600
net2599
net2598
net2597
net2596
net2595
net2594
net2593
net2592
net2591
net2590
net2589
net2588
net2587
net2586
net2585
net2584
net2583
net2582
net2581
net2580
net2579
net2578
net2577
net2576
net2575
net2574
net2573
net2572
net2571
net2570
net2569
net2568
net2567
net2566
net2565
net2564
net2563
net2562
net2561
net2560
net2559
net2558
net2557
net2556
net2555
net2554
net2553
net2552
net2551
net2550
net2549
net2548
net2547
net2546
net2545
net2544
net2543
net2542
net2541
net2540
net2539
net2538
net2537
net2536
net2535
net2534
net2533
net2532
net2531
net2530
net2529
net2528
net2527
net2526
net2525
net2524
net2523
net2522
net2521
net2520
net2519
net2518
net2517
net2516
net2515
net2514
net2513
net2512
net2511
net2510
net2509
net2508
net2507
net2506
net2505
net2504
net2503
net2502
net2501
net2500
net2499
net2498
net2497
net2496
net2495
net2494
net2493
net2492
net2491
net2490
net2489
net2488
net2487
net2486
net2485
net2484
net2483
net2482
net2481
net2480
net2479
net2478
net2477
net2476
net2475
net2474
net2473
net2472
net2471
net2470
net2469
net2468
net2467
net2466
net2465
net2464
net2463
net2462
net2461
net2460
net2459
net2458
net2457
net2456
net2455
net2454
net2453
net2452
net2451
net2450
net2449
net2448
net2447
net2446
net2445
net2444
net2443
net2441
net2440
net2439
net2438
net2437
net2436
net2435
net2434
net2433
net2432
net2431
net2430
net2429
net2428
net2427
net2426
net2425
net2424
net2423
net2422
net2421
net2420
net2419
net2418
net2417
net2416
net2415
net2414
net2413
net2412
net2411
net2410
net2409
net2408
net2407
net2406
net2405
net2404
net2403
net2402
net2401
net2400
net2399
net2398
net2397
net2396
net2395
net2394
net2393
net2392
net2391
net2390
net2389
net2388
net2387
net2386
net2385
net2384
net2383
net2382
net2381
net2380
net2379
net2378
net2377
net2376
net2375
net2374
net2373
net2372
net2371
net2370
net2369
net2368
net2367
net2366
net2365
net2364
net2363
net2362
net2361
net2360
net2359
net2358
net2357
net2356
net2355
net2354
net2353
net2352
net2351
net2350
net2349
net2348
net2347
net2346
net2345
net2344
net2343
net2342
net2341
net2340
net2339
net2338
net2337
net2336
net2335
net2334
net2333
net2332
net2331
net2330
net2329
net2328
net2327
net2326
net2325
net2324
net2323
net2322
net2321
net2320
net2319
net2318
net2317
net2316
net2315
net2314
net2313
net2312
net2311
net2310
net2309
net2308
net2307
net2306
net2305
net2303
net2302
net2301
net2300
net2299
net2298
net2297
net2296
net2295
net2294
net2293
net2292
net2291
net2290
net2289
net2288
net2287
net2286
net2285
net2284
net2283
net2282
net2281
net2280
net2279
net2278
net2277
net2276
net2275
net2274
net2273
net2272
net2271
net2270
net2269
net2268
net2267
net2266
net2265
net2264
net2263
net2262
net2261
net2260
net2259
net2258
net2257
net2256
net2255
net2254
net2253
net2252
net2251
net2250
net2249
net2248
net2247
net2246
net2245
net2244
net2243
net2242
net2241
net2240
net2239
net2238
net2237
net2236
net2235
net2234
net2233
net2232
net2231
net2230
net2229
net2228
net2227
net2226
net2225
net2224
net2223
net2222
net2221
net2220
net2219
net2218
net2217
net2216
net2215
net2214
net2213
net2212
net2211
net2210
net2209
net2208
net2207
net2206
net2205
net2204
net2203
net2202
net2201
net2200
net2199
net2198
net2197
net2196
net2195
net2194
net2193
net2192
net2191
net2190
net2189
net2188
net2187
net2186
net2185
net2184
net2183
net2182
net2181
net2180
net2179
net2178
net2177
net2176
net2175
net2174
net2173
net2172
net2171
net2170
net2169
net2168
net2167
net2166
net2165
net2164
net2163
net2162
net2161
net2160
net2159
net2158
net2157
net2156
net2155
net2154
net2153
net2152
net2151
net2150
net2149
net2148
net2147
net2146
net2145
net2144
net2143
net2141
net2140
net2139
net2138
net2137
net2136
net2135
net2134
net2133
net2132
net2131
net2130
net2129
net2128
net2127
net2126
net2125
net2124
net2123
net2122
net2121
net2120
net2119
net2118
net2117
net2116
net2115
net2114
net2113
net2112
net2111
net2110
net2109
net2108
net2107
net2106
net2105
net2104
net2103
net2102
net2101
net2100
net2099
net2098
net2097
net2096
net2095
net2094
net2093
net2092
net2091
net2090
net2089
net2088
net2087
net2086
net2085
net2084
net2083
net2082
net2081
net2080
net2079
net2078
net2077
net2076
net2075
net2074
net2073
net2072
net2071
net2070
net2069
net2068
net2067
net2066
net2065
net2064
net2063
net2062
net2061
net2060
net2059
net2058
net2057
net2056
net2055
net2054
net2053
net2052
net2051
net2050
net2049
net2048
net2047
net2046
net2045
net2044
net2043
net2042
net2041
net2040
net2039
net2038
net2037
net2036
net2035
net2034
net2033
net2032
net2031
net2030
net2029
net2028
net2027
net2026
net2025
net2024
net2023
net2022
net2021
net2020
net2019
net2018
net2017
net2016
net2015
net2014
net2013
net2012
net2011
net2010
net2009
net2008
net2007
net2006
net2005
net2004
net2003
net2002
net2001
net2000
net1999
net1998
net1997
net1996
net1995
net1994
net1993
net1992
net1991
net1990
net1989
net1988
net1987
net1986
net1985
net1984
net1983
net1982
net1981
net1980
net1979
net1978
net1977
net1976
net1975
net1974
net1973
net1972
net1971
net1970
net1969
net1968
net1967
net1966
net1965
net1964
net1963
net1962
net1961
net1960
net1959
net1958
net1957
net1956
net1955
net1954
net1953
net1952
net1951
net1950
net1949
net1948
net1947
net1946
net1945
net1944
net1943
net1942
net1941
net1940
net1939
net1938
net1937
net1936
net1935
net1934
net1933
net1932
net1931
net1930
net1929
net1928
net1927
net1926
net1925
net1924
net1923
net1922
net1921
net1920
net1919
net1918
net1917
net1916
net1915
net1914
net1913
net1912
net1911
net1910
net1909
net1908
net1907
net1906
net1905
net1904
net1903
net1902
net1901
net1900
net1899
net1898
net1897
net1896
net1895
net1894
net1893
net1892
net1891
net1890
net1889
net1888
net1887
net1886
net1885
net1884
net1883
net1882
net1881
net1880
net1879
net1878
net1877
net1876
net1875
net1874
net1873
net1872
net1871
net1870
net1869
net1868
net1867
net1866
net1865
net1864
net1863
net1862
net1861
net1860
net1859
net1858
net1857
net1856
net1855
net1854
net1853
net1852
net1851
net1850
net1849
net1848
net1847
net1846
net1845
net1844
net1843
net1842
net1841
net1840
net1839
net1838
net1837
net1836
net1835
net1834
net1833
net1832
net1831
net1830
net1829
net1828
net1827
net1826
net1825
net1824
net1823
net1822
net1821
net1820
net1819
net1818
net1817
net1816
net1815
net1814
net1813
net1812
net1811
net1810
net1809
net1808
net1807
net1806
net1805
net1804
net1803
net1802
net1801
net1800
net1799
net1798
net1797
net1796
net1795
net1794
net1792
net1791
net1790
net1789
net1788
net1787
net1786
net1785
net1784
net1783
net1782
net1781
net1780
net1779
net1778
net1777
net1776
net1775
net1774
net1773
net1772
net1771
net1770
net1769
net1768
net1767
net1766
net1765
net1764
net1763
net1762
net1761
net1760
net1759
net1758
net1757
net1756
net1755
net1754
net1753
net1752
net1751
net1750
net1749
net1748
net1747
net1746
net1745
net1744
net1743
net1742
net1741
net1740
net1739
net1738
net1737
net1736
net1735
net1734
net1733
net1732
net1731
net1730
net1729
net1728
net1727
net1726
net1725
net1724
net1723
net1722
net1721
net1720
net1719
net1718
net1717
net1716
net1715
net1714
net1713
net1712
net1711
net1710
net1709
net1708
net1707
net1706
net1705
net1704
net1703
net1702
net1701
net1700
net1699
net1698
net1697
net1696
net1695
net1694
net1693
net1692
net1691
net1690
net1689
net1688
net1687
net1686
net1685
net1684
net1683
net1682
net1681
net1680
net1679
net1678
net1677
net1676
net1675
net1674
net1673
net1672
net1671
net1670
net1669
net1668
net1667
net1666
net1665
net1664
net1663
net1662
net1661
net1660
net1659
net1657
net1656
net1655
net1654
net1653
net1652
net1651
net1650
net1649
net1648
net1647
net1646
net1645
net1644
net1643
net1642
net1641
net1640
net1639
net1638
net1637
net1636
net1635
net1634
net1633
net1632
net1631
net1630
net1629
net1628
net1627
net1626
net1625
net1624
net1623
net1622
net1621
net1620
net1619
net1618
net1617
net1616
net1615
net1614
net1613
net1612
net1611
net1610
net1609
net1608
net1607
net1606
net1605
net1604
net1603
net1602
net1601
net1600
net1599
net1598
net1597
net1596
net1595
net1594
net1593
net1592
net1591
net1590
net1589
net1588
net1587
net1586
net1585
net1584
net1583
net1582
net1581
net1580
net1579
net1578
net1577
net1576
net1575
net1574
net1573
net1572
net1571
net1570
net1569
net1568
net1567
net1566
net1565
net1564
net1563
net1562
net1561
net1560
net1559
net1558
net1557
net1556
net1555
net1554
net1553
net1552
net1551
net1550
net1549
net1548
net1547
net1546
net1545
net1544
net1543
net1542
net1541
net1540
net1539
net1538
net1537
net1536
net1535
net1534
net1533
net1532
net1531
net1529
net1528
net1527
net1526
net1525
net1524
net1523
net1522
net1521
net1520
net1519
net1518
net1517
net1516
net1515
net1514
net1513
net1512
net1511
net1510
net1509
net1508
net1507
net1506
net1505
net1504
net1503
net1502
net1501
net1500
net1499
net1498
net1497
net1496
net1495
net1494
net1493
net1492
net1491
net1490
net1489
net1488
net1487
net1486
net1485
net1484
net1483
net1482
net1481
net1480
net1479
net1478
net1477
net1476
net1475
net1474
net1473
net1472
net1471
net1470
net1469
net1468
net1467
net1466
net1465
net1464
net1463
net1462
net1461
net1460
net1459
net1458
net1457
net1456
net1455
net1454
net1453
net1452
net1451
net1450
net1449
net1448
net1447
net1446
net1445
net1444
net1443
net1442
net1441
net1440
net1439
net1438
net1437
net1436
net1435
net1434
net1433
net1432
net1431
net1430
net1429
net1428
net1427
net1426
net1425
net1424
net1423
net1422
net1421
net1420
net1419
net1418
net1417
net1416
net1415
net1414
net1413
net1412
net1411
net1410
net1409
net1408
net1407
net1406
net1405
net1404
net1403
net1402
net1401
net1400
net1399
net1398
net1397
net1396
net1395
net1394
net1393
net1392
net1391
net1390
net1389
net1388
net1387
net1386
net1385
net1384
net1383
net1382
net1381
net1380
net1379
net1378
net1377
net1376
net1375
net1374
net1373
net1372
net1371
net1370
net1369
net1368
net1367
net1366
net1365
net1364
net1363
net1362
net1361
net1360
net1359
net1358
net1357
net1356
net1355
net1354
net1353
net1352
net1351
net1350
net1349
net1348
net1347
net1346
net1345
net1344
net1343
net1342
net1341
net1340
net1339
net1338
net1337
net1336
net1335
net1334
net1333
net1332
net1331
net1330
net1329
net1328
net1327
net1326
net1325
net1324
net1323
net1322
net1321
net1320
net1319
net1318
net1317
net1316
net1315
net1314
net1313
net1312
net1311
net1310
net1309
net1308
net1307
net1306
net1305
net1304
net1303
net1302
net1301
net1300
net1299
net1298
net1297
net1296
net1295
net1294
net1293
net1292
net1291
net1290
net1289
net1288
net1287
net1286
net1285
net1284
net1283
net1282
net1281
net1280
net1279
net1278
net1277
net1276
net1275
net1274
net1273
net1272
net1271
net1270
net1269
net1268
net1267
net1266
net1265
net1264
net1263
net1262
net1261
net1260
net1259
net1258
net1257
net1256
net1255
net1254
net1253
net1252
net1251
net1250
net1249
net1248
net1247
net1246
net1245
net1244
net1243
net1242
net1241
net1240
net1239
net1238
net1237
net1236
net1235
net1234
net1233
net1232
net1231
net1230
net1229
net1228
net1227
net1226
net1225
net1224
net1223
net1222
net1221
net1220
net1219
net1218
net1217
net1216
net1215
net1214
net1213
net1212
net1211
net1210
net1209
net1208
net1207
net1206
net1205
net1204
net1203
net1202
net1201
net1200
net1199
net1198
net1197
net1196
net1195
net1194
net1193
net1192
net1191
net1190
net1189
net1188
net1187
net1186
net1185
net1184
net1183
net1182
net1181
net1180
net1179
net1178
net1177
net1176
net1175
net1174
net1173
net1172
net1171
net1170
net1169
net1168
net1167
net1166
net1165
net1164
net1163
net1162
net1161
net1160
net1159
net1158
net1157
net1156
net1155
net1154
net1153
net1152
net1151
net1150
net1149
net1148
net1147
net1146
net1145
net1144
net1143
net1142
net1141
net1140
net1139
net1138
net1137
net1136
net1135
net1134
net1133
net1132
net1131
net1130
net1129
net1128
net1127
net1126
net1125
net1124
net1123
net1122
net1121
net1120
net1119
net1118
net1117
net1116
net1115
net1114
net1113
net1112
net1111
net1110
net1109
net1108
net1107
net1106
net1105
net1104
net1103
net1102
net1101
net1100
net1099
net1098
net1097
net1096
net1095
net1094
net1093
net1092
net1091
net1090
net1089
net1088
net1087
net1086
net1085
net1084
net1083
net1082
net1081
net1080
net1079
net1078
net1077
net1076
net1075
net1074
net1073
net1072
net1071
net1070
net1069
net1068
net1067
net1066
net1065
net1064
net1063
net1062
net1061
net1060
net1059
net1058
net1057
net1056
net1055
net1054
net1053
net1052
net1051
net1050
net1049
net1048
net1047
net1046
net1045
net1044
net1043
net1042
net1041
net1040
net1039
net1038
net1037
net1036
net1035
net1034
net1033
net1032
net1031
net1030
net1029
net1028
net1027
net1026
net1025
net1024
net1023
net1022
net1021
net1020
net1019
net1018
net1017
net1016
net1015
net1014
net1013
net1012
net1011
net1010
net1009
net1008
net1007
net1006
net1005
net1004
net1003
net1002
net1001
net1000
net999
net998
net997
net996
net995
net994
net993
net992
net991
net990
net989
net988
net987
net986
net985
net984
net983
net982
net981
net980
net979
net978
net977
net976
net975
net974
net973
net972
net971
net970
net969
net968
net967
net966
net965
net964
net963
net962
net961
net960
net959
net958
net957
net956
net955
net954
net953
net952
net951
net950
net949
net948
net947
net946
net945
net944
net943
net942
net941
net940
net939
net938
net937
net936
net935
net934
net933
net932
net931
net930
net928
net927
net926
net925
net924
net923
net922
net921
net920
net919
net918
net917
net916
net915
net914
net913
net912
net911
net910
net909
net908
net907
net906
net905
net904
net903
net902
net901
net900
net899
net898
net897
net896
net895
net894
net893
net892
net891
net890
net889
net888
net887
net886
net885
net884
net883
net882
net881
net880
net879
net878
net877
net876
net875
net874
net873
net872
net871
net870
net869
net868
net867
net866
net865
net864
net863
net862
net861
net860
net859
net858
net857
net856
net855
net854
net853
net852
net851
net850
net849
net848
net847
net846
net845
net844
net843
net842
net841
net840
net839
net838
net837
net836
net835
net834
net833
net832
net831
net829
net828
net827
net826
net825
net824
net823
net822
net821
net820
net819
net818
net817
net816
net815
net814
net813
net812
net811
net810
net809
net808
net807
net806
net805
net804
net803
net802
net801
net800
net799
net798
net797
net795
net794
net793
net792
net791
net790
net789
net788
net787
net786
net785
net784
net783
net782
net781
net780
net779
net778
net777
net776
net775
net774
net773
net772
net771
net770
net769
net768
net767
net766
net765
net764
net763
net762
net761
net760
net759
net758
net757
net756
net755
net754
net753
net752
net751
net750
net749
net748
net747
net746
net745
net744
net743
net742
net741
net740
net739
net738
net737
net735
net734
net733
net732
net731
net730
net729
net728
net727
net726
net725
net724
net723
net722
net721
net720
net719
net718
net717
net716
net715
net714
net713
net712
net711
net710
net709
net708
net707
net706
net705
net704
net703
net702
net701
net700
net699
net698
net697
net696
net695
net694
net693
net692
net691
net690
net689
net688
net687
net686
net685
net684
net683
net682
net681
net680
net679
net678
net677
net676
net675
net674
net673
net672
net671
net670
net669
net668
net667
net666
net665
net664
net663
net662
net661
net660
net659
net658
net657
net656
net655
net654
net653
net652
net651
net650
net649
net648
net647
net646
net645
net644
net643
net642
net641
net640
net639
net638
net637
net636
net635
net634
net633
net632
net631
net630
net629
net628
net627
net626
net625
net624
net623
net621
net620
net619
net618
net617
net616
net615
net614
net613
net612
net611
net610
net609
net608
net607
net606
net605
net604
net603
net602
net601
net600
net599
net598
net597
net596
net595
net594
net593
net592
net591
net590
net589
net588
net587
net586
net585
net584
net583
net582
net581
net580
net579
net578
net577
net576
net575
net574
net573
net572
net571
net570
net569
net568
net567
net566
net565
net564
net563
net562
net561
net560
net559
net558
net557
net556
net555
net554
net553
net552
net551
net550
net549
net548
net547
net546
net545
net544
net543
net542
net541
net540
net539
net538
net537
net536
net535
net534
net533
net532
net531
net530
net529
net528
net527
net526
net525
net524
net523
net522
net521
net520
net519
net518
net517
net516
net515
net514
net513
net512
net511
net510
net509
net508
net507
net506
net505
net504
net503
net502
net501
net500
net499
net498
net497
net496
net495
net494
net493
net492
net491
net490
net489
net488
net487
net486
net485
net484
net483
net482
net481
net480
net479
net478
net477
net476
net475
net474
net473
net472
net471
net470
net469
net468
net467
net466
net465
net464
net463
net462
net461
net460
net459
net458
net457
net456
net455
net454
net453
net452
net451
net450
net449
net448
net447
net445
net444
net443
net442
net441
net440
net439
net438
net437
net436
net435
net434
net433
net432
net431
net430
net429
net428
net427
net426
net425
net424
net423
net422
net421
net420
net419
net418
net417
net416
net415
net414
net413
net412
net411
net410
net409
net408
net407
net406
net404
net403
net402
net401
net400
net399
net398
net397
net396
net395
net394
net393
net392
net391
net390
net389
net388
net387
net386
net385
net384
net383
net382
net381
net380
net379
net378
net377
net376
net375
net374
net373
net372
net371
net370
net369
net368
net367
net366
net365
net364
net363
net362
net361
net360
net359
net358
net357
net356
net355
net354
net353
net352
net351
net350
net349
net348
net347
net346
net345
net344
net343
net342
net341
net340
net339
net338
net337
net336
net335
net334
net333
net332
net331
net330
net329
net328
net327
net326
net325
net324
net323
net322
net321
net320
net319
net318
net317
net316
net315
net314
net313
net312
net311
net310
net309
net308
net307
net306
net305
net304
net303
net302
net301
net300
net299
net298
net297
net296
net295
net294
net293
net292
net291
net290
net289
net288
net287
net286
net285
net284
net283
net282
net281
net280
net279
net278
net277
net276
net275
net274
net273
net272
net271
net270
net269
net268
net267
net266
net265
net264
net263
net262
net261
net260
net259
net258
net257
net256
net255
net254
net253
net252
net251
net250
net249
net248
net247
net246
net245
net244
net243
net242
net241
net240
net239
net238
net237
net236
net235
net234
net233
net232
net231
net230
net229
net228
net227
net226
net225
net224
net223
net222
net221
net220
net219
net218
net217
net216
net215
net214
net213
net212
net211
net210
net209
net208
net207
net206
net205
net204
net203
net202
net201
net200
net199
net198
net197
net196
net195
net194
net193
net192
net191
net190
net189
net188
net187
net186
net185
net184
net183
net182
net181
net180
net179
net178
net177
net176
net175
net174
net173
net172
net171
net170
net169
net168
net167
net166
net165
net164
net163
net162
net161
net160
net159
net158
net157
net156
net155
net154
net153
net152
net151
net150
net149
net147
net146
net145
net144
net143
net142
net141
net140
net139
net138
net137
net136
net135
net134
net133
net132
net131
net130
net129
net128
net127
net126
net125
net124
net123
net122
net121
net120
net119
net118
net117
net116
net115
net114
net113
net112
net111
net110
net109
net108
net107
net106
net105
net104
net103
net102
net101
net100
net99
net98
net97
net96
net95
net94
net93
net92
net91
net90
net89
net88
net87
net86
net85
net84
net83
net82
net81
net80
net79
net78
net77
net76
net75
net74
net73
net72
net71
net70
net69
net68
net67
net66
net65
net64
net63
net62
net61
net60
net59
net58
net57
net56
net55
net54
net53
net52
net51
net50
net49
net48
net47
net46
net45
net44
net43
net42
net41
net40
net39
net38
net37
net36
net35
net34
net33
net32
net31
net30
net29
net28
net27
net26
net25
net24
net23
net22
net21
net20
net19
net18
net17
net16
net15
net14
net13
net12
net11
net10
net9
net8
net7
net5
net4
net3
net2
net1
net0
XOR2XL
--pins(5)
Y
use :  
dir : o
shape : 
(2582,558):(2704,1590) : 0
(2524,558):(2582,720) : 0
(2564,1146):(2582,1254) : 0
(2524,1428):(2582,1590) : 0
B
use :  
dir : i
shape : 
(700,1140):(758,1250) : 0
(578,1140):(700,1522) : 0
(464,1412):(578,1522) : 0
A
use :  
dir : i
shape : 
(1002,1114):(1084,1276) : 0
(880,878):(1002,1276) : 0
(814,878):(880,992) : 0
(464,884):(814,992) : 0
(446,866):(464,992) : 0
(324,776):(446,992) : 0
VSS
use : g
dir : b
shape : 
(2408,-160):(2800,160) : 0
(2228,-160):(2408,244) : 0
(650,-160):(2228,160) : 0
(470,-160):(650,244) : 0
(0,-160):(470,160) : 0
VDD
use : p
dir : b
shape : 
(2408,2240):(2800,2560) : 0
(2228,2156):(2408,2560) : 0
(610,2240):(2228,2560) : 0
(430,2156):(610,2560) : 0
(0,2240):(430,2560) : 0
XOR2X4
--pins(5)
Y
use :  
dir : o
shape : 
(5450,672):(5572,2066) : 0
(5358,672):(5450,834) : 0
(5368,1400):(5450,2066) : 0
(5358,1452):(5368,1678) : 0
B
use :  
dir : i
shape : 
(590,1000):(796,1162) : 0
(468,1000):(590,1254) : 0
(294,1000):(468,1162) : 0
A
use :  
dir : i
shape : 
(3998,1100):(4120,1254) : 0
(3776,1100):(3998,1210) : 0
(3594,1048):(3776,1210) : 0
VSS
use : g
dir : b
shape : 
(5904,-160):(6000,160) : 0
(5722,-160):(5904,244) : 0
(5176,-160):(5722,160) : 0
(4994,-160):(5176,244) : 0
(4374,-160):(4994,160) : 0
(4192,-160):(4374,244) : 0
(1668,-160):(4192,160) : 0
(1486,-160):(1668,244) : 0
(962,-160):(1486,160) : 0
(780,-160):(962,456) : 0
(278,-160):(780,160) : 0
(96,-160):(278,456) : 0
(0,-160):(96,160) : 0
VDD
use : p
dir : b
shape : 
(5904,2240):(6000,2560) : 0
(5722,2156):(5904,2560) : 0
(5176,2240):(5722,2560) : 0
(4994,2156):(5176,2560) : 0
(4406,2240):(4994,2560) : 0
(4224,2156):(4406,2560) : 0
(1668,2240):(4224,2560) : 0
(1486,2156):(1668,2560) : 0
(962,2240):(1486,2560) : 0
(780,1978):(962,2560) : 0
(278,2240):(780,2560) : 0
(96,1978):(278,2560) : 0
(0,2240):(96,2560) : 0
XOR2X2
--pins(5)
Y
use :  
dir : o
shape : 
(3370,342):(3496,1996) : 0
(3310,342):(3370,790) : 0
(3310,1386):(3370,1996) : 0
B
use :  
dir : i
shape : 
(736,1128):(922,1388) : 0
(652,1278):(736,1388) : 0
(526,1278):(652,1526) : 0
(478,1412):(526,1526) : 0
A
use :  
dir : i
shape : 
(1738,998):(1862,1170) : 0
(1372,1060):(1738,1170) : 0
(1274,1060):(1372,1260) : 0
(1148,908):(1274,1260) : 0
(458,908):(1148,1016) : 0
(332,908):(458,1110) : 0
VSS
use : g
dir : b
shape : 
(3066,-160):(3600,160) : 0
(2880,-160):(3066,244) : 0
(1440,-160):(2880,160) : 0
(1254,-160):(1440,244) : 0
(610,-160):(1254,160) : 0
(426,-160):(610,244) : 0
(0,-160):(426,160) : 0
VDD
use : p
dir : b
shape : 
(3060,2240):(3600,2560) : 0
(2874,2156):(3060,2560) : 0
(1396,2240):(2874,2560) : 0
(1210,1810):(1396,2560) : 0
(610,2240):(1210,2560) : 0
(426,1810):(610,2560) : 0
(0,2240):(426,2560) : 0
XOR2X1
--pins(5)
Y
use :  
dir : o
shape : 
(2582,558):(2704,1576) : 0
(2524,558):(2582,720) : 0
(2564,1146):(2582,1576) : 0
(2524,1414):(2564,1576) : 0
B
use :  
dir : i
shape : 
(700,1140):(758,1250) : 0
(578,1140):(700,1522) : 0
(464,1412):(578,1522) : 0
A
use :  
dir : i
shape : 
(1002,1114):(1084,1276) : 0
(880,878):(1002,1276) : 0
(814,878):(880,992) : 0
(464,884):(814,992) : 0
(446,866):(464,992) : 0
(324,776):(446,992) : 0
VSS
use : g
dir : b
shape : 
(2408,-160):(2800,160) : 0
(2228,-160):(2408,244) : 0
(650,-160):(2228,160) : 0
(470,-160):(650,244) : 0
(0,-160):(470,160) : 0
VDD
use : p
dir : b
shape : 
(2408,2240):(2800,2560) : 0
(2228,2156):(2408,2560) : 0
(610,2240):(2228,2560) : 0
(430,2156):(610,2560) : 0
(0,2240):(430,2560) : 0
XNOR2X4
--pins(5)
Y
use :  
dir : o
shape : 
(5450,672):(5572,2066) : 0
(5358,672):(5450,834) : 0
(5368,1400):(5450,2066) : 0
(5358,1452):(5368,1614) : 0
B
use :  
dir : i
shape : 
(590,1000):(796,1162) : 0
(468,1000):(590,1254) : 0
(294,1000):(468,1162) : 0
A
use :  
dir : i
shape : 
(1714,1034):(1894,1196) : 0
(1526,1034):(1714,1254) : 0
VSS
use : g
dir : b
shape : 
(5904,-160):(6000,160) : 0
(5722,-160):(5904,244) : 0
(5176,-160):(5722,160) : 0
(4994,-160):(5176,244) : 0
(4374,-160):(4994,160) : 0
(4192,-160):(4374,244) : 0
(1668,-160):(4192,160) : 0
(1486,-160):(1668,244) : 0
(962,-160):(1486,160) : 0
(780,-160):(962,456) : 0
(278,-160):(780,160) : 0
(96,-160):(278,456) : 0
(0,-160):(96,160) : 0
VDD
use : p
dir : b
shape : 
(5904,2240):(6000,2560) : 0
(5722,2156):(5904,2560) : 0
(5176,2240):(5722,2560) : 0
(4994,2156):(5176,2560) : 0
(4406,2240):(4994,2560) : 0
(4224,2156):(4406,2560) : 0
(1668,2240):(4224,2560) : 0
(1486,2156):(1668,2560) : 0
(962,2240):(1486,2560) : 0
(780,1978):(962,2560) : 0
(278,2240):(780,2560) : 0
(96,1978):(278,2560) : 0
(0,2240):(96,2560) : 0
XNOR2X2
--pins(5)
Y
use :  
dir : o
shape : 
(3896,342):(3900,790) : 0
(3768,342):(3896,1996) : 0
(3714,342):(3768,790) : 0
(3708,1386):(3768,1996) : 0
B
use :  
dir : i
shape : 
(980,1128):(1042,1290) : 0
(854,1128):(980,1388) : 0
(804,1254):(854,1388) : 0
(658,1278):(804,1388) : 0
(532,1278):(658,1526) : 0
(482,1412):(532,1526) : 0
A
use :  
dir : i
shape : 
(2118,936):(2246,1170) : 0
(1750,1060):(2118,1170) : 0
(1622,1060):(1750,1260) : 0
(1336,1150):(1622,1260) : 0
(1294,1146):(1336,1260) : 0
(1168,908):(1294,1260) : 0
(462,908):(1168,1016) : 0
(336,908):(462,1110) : 0
VSS
use : g
dir : b
shape : 
(3482,-160):(4000,160) : 0
(3294,-160):(3482,244) : 0
(1620,-160):(3294,160) : 0
(1432,-160):(1620,244) : 0
(772,-160):(1432,160) : 0
(584,-160):(772,244) : 0
(0,-160):(584,160) : 0
VDD
use : p
dir : b
shape : 
(3454,2240):(4000,2560) : 0
(3268,2156):(3454,2560) : 0
(1576,2240):(3268,2560) : 0
(1388,1810):(1576,2560) : 0
(760,2240):(1388,2560) : 0
(574,1810):(760,2560) : 0
(0,2240):(574,2560) : 0
XNOR2X1
--pins(5)
Y
use :  
dir : o
shape : 
(2582,558):(2704,1576) : 0
(2524,558):(2582,720) : 0
(2564,1146):(2582,1576) : 0
(2524,1414):(2564,1576) : 0
B
use :  
dir : i
shape : 
(700,1110):(758,1272) : 0
(578,1110):(700,1522) : 0
(464,1412):(578,1522) : 0
A
use :  
dir : i
shape : 
(1002,1114):(1084,1276) : 0
(880,878):(1002,1276) : 0
(814,878):(880,992) : 0
(464,884):(814,992) : 0
(446,878):(464,992) : 0
(324,776):(446,992) : 0
VSS
use : g
dir : b
shape : 
(2408,-160):(2800,160) : 0
(2228,-160):(2408,244) : 0
(650,-160):(2228,160) : 0
(470,-160):(650,244) : 0
(0,-160):(470,160) : 0
VDD
use : p
dir : b
shape : 
(2408,2240):(2800,2560) : 0
(2228,2156):(2408,2560) : 0
(636,2240):(2228,2560) : 0
(456,2156):(636,2560) : 0
(0,2240):(456,2560) : 0
SEDFFXL
--pins(9)
SI
use :  
dir : i
shape : 
(1462,1066):(1746,1266) : 0
SE
use :  
dir : i
shape : 
(664,1086):(932,1300) : 0
QN
use :  
dir : o
shape : 
(9166,758):(9286,1648) : 0
(9036,758):(9166,866) : 0
(9010,1486):(9166,1648) : 0
(8856,642):(9036,866) : 0
Q
use :  
dir : o
shape : 
(8600,426):(8722,1784) : 0
(8468,426):(8600,536) : 0
(8590,1674):(8600,1784) : 0
(8468,1674):(8590,1800) : 0
(8348,334):(8468,536) : 0
(8408,1690):(8468,1800) : 0
(8286,1690):(8408,2012) : 0
(8168,324):(8348,536) : 0
(8228,1850):(8286,2012) : 0
E
use :  
dir : i
shape : 
(462,1678):(582,1820) : 0
(372,1710):(462,1820) : 0
(250,1710):(372,1962) : 0
(192,1800):(250,1962) : 0
D
use :  
dir : i
shape : 
(2110,1048):(2364,1254) : 0
CK
use : c
dir : i
shape : 
(4900,866):(5148,1084) : 0
VSS
use : g
dir : b
shape : 
(8992,-160):(9400,160) : 0
(8812,-160):(8992,244) : 0
(7908,-160):(8812,160) : 0
(7786,-160):(7908,716) : 0
(6460,-160):(7786,160) : 0
(6280,-160):(6460,436) : 0
(5530,-160):(6280,160) : 0
(5352,-160):(5530,384) : 0
(1714,-160):(5352,160) : 0
(1594,-160):(1714,398) : 0
(348,-160):(1594,160) : 0
(168,-160):(348,244) : 0
(0,-160):(168,160) : 0
VDD
use : p
dir : b
shape : 
(9072,2240):(9400,2560) : 0
(8864,2156):(9072,2560) : 0
(8004,2226):(8864,2560) : 0
(7826,1650):(8004,2560) : 0
(6592,2240):(7826,2560) : 0
(6096,2156):(6592,2560) : 0
(5518,2240):(6096,2560) : 0
(4726,2156):(5518,2560) : 0
(1556,2240):(4726,2560) : 0
(1376,1926):(1556,2560) : 0
(744,2240):(1376,2560) : 0
(564,1972):(744,2560) : 0
(0,2240):(564,2560) : 0
SEDFFX4
--pins(9)
SI
use :  
dir : i
shape : 
(1770,1058):(2084,1266) : 0
SE
use : �
dir : i
shape : 
(686,1086):(1048,1254) : 0
QN
use : �
dir : o
shape : 
(11428,664):(11732,826) : 0
(11418,1380):(11646,1542) : 0
(11418,600):(11428,1266) : 0
(11238,600):(11418,1542) : 0
(11228,600):(11238,1266) : 0
Q
use : 
dir : o
shape : 
(11070,600):(11080,1266) : 0
(10890,600):(11070,1542) : 0
(10880,600):(10890,1266) : 0
(10790,1380):(10890,1542) : 0
(10878,662):(10880,824) : 0
E
use : z
dir : i
shape : 
(530,1678):(584,1788) : 0
(410,1678):(530,1910) : 0
(390,1800):(410,1910) : 0
(212,1800):(390,1962) : 0
D
use : z
dir : i
shape : 
(2614,1146):(2676,1254) : 0
(2406,1146):(2614,1388) : 0
CK
use : c
dir : i
shape : 
(5144,866):(5504,1058) : 0
VSS
use : g
dir : b
shape : 
(12104,-160):(12200,160) : 0
(11926,-160):(12104,494) : 0
(11394,-160):(11926,160) : 0
(11216,-160):(11394,442) : 0
(10716,-160):(11216,160) : 0
(10536,-160):(10716,424) : 0
(9966,-160):(10536,160) : 0
(9786,-160):(9966,770) : 0
(8510,-160):(9786,160) : 0
(8332,-160):(8510,244) : 0
(7138,-160):(8332,160) : 0
(6958,-160):(7138,450) : 0
(5884,-160):(6958,160) : 0
(5704,-160):(5884,446) : 0
(1804,-160):(5704,160) : 0
(1624,-160):(1804,432) : 0
(338,-160):(1624,160) : 0
(158,-160):(338,244) : 0
(0,-160):(158,160) : 0
VDD
use : p
dir : b
shape : 
(12004,2240):(12200,2560) : 0
(11826,1930):(12004,2560) : 0
(11308,2240):(11826,2560) : 0
(11128,1978):(11308,2560) : 0
(10632,2240):(11128,2560) : 0
(10452,1978):(10632,2560) : 0
(9850,2240):(10452,2560) : 0
(9622,2156):(9850,2560) : 0
(8356,2240):(9622,2560) : 0
(8176,2156):(8356,2560) : 0
(6848,2240):(8176,2560) : 0
(6668,2156):(6848,2560) : 0
(5654,2240):(6668,2560) : 0
(5474,2156):(5654,2560) : 0
(4964,2240):(5474,2560) : 0
(4784,2156):(4964,2560) : 0
(1728,2240):(4784,2560) : 0
(1548,1882):(1728,2560) : 0
(924,2240):(1548,2560) : 0
(744,1840):(924,2560) : 0
(0,2240):(744,2560) : 0
SEDFFX2
--pins(9)
SI
use :  
dir : i
shape : 
(1482,1066):(1750,1266) : 0
SE
use : �
dir : i
shape : 
(746,1040):(996,1284) : 0
QN
use :  
dir : o
shape : 
(10184,612):(10306,1920) : 0
(10166,612):(10184,812) : 0
(10126,1472):(10184,1920) : 0
(10106,650):(10166,812) : 0
Q
use : 
dir : o
shape : 
(9594,650):(9610,878) : 0
(9580,612):(9594,878) : 0
(9518,612):(9580,1412) : 0
(9460,612):(9518,1524) : 0
(9434,650):(9460,878) : 0
(9396,1210):(9460,1524) : 0
(9430,650):(9434,812) : 0
E
use :  
dir : i
shape : 
(486,1678):(580,1788) : 0
(394,1678):(486,1910) : 0
(366,1678):(394,1962) : 0
(216,1800):(366,1962) : 0
D
use :  
dir : i
shape : 
(2056,1074):(2354,1266) : 0
CK
use : c
dir : i
shape : 
(4926,866):(5144,1128) : 0
VSS
use : g
dir : b
shape : 
(9948,-160):(10400,160) : 0
(9770,-160):(9948,442) : 0
(8896,-160):(9770,160) : 0
(8716,-160):(8896,636) : 0
(7844,-160):(8716,160) : 0
(8714,534):(8716,634) : 0
(7666,-160):(7844,474) : 0
(6456,-160):(7666,160) : 0
(6276,-160):(6456,380) : 0
(5520,-160):(6276,160) : 0
(5342,-160):(5520,398) : 0
(1792,-160):(5342,160) : 0
(1612,-160):(1792,358) : 0
(336,-160):(1612,160) : 0
(158,-160):(336,244) : 0
(0,-160):(158,160) : 0
VDD
use : p
dir : b
shape : 
(9928,2240):(10400,2560) : 0
(9748,1970):(9928,2560) : 0
(8780,2234):(9748,2560) : 0
(7992,2156):(8780,2560) : 0
(6542,2240):(7992,2560) : 0
(6006,2156):(6542,2560) : 0
(5312,2240):(6006,2560) : 0
(4640,2156):(5312,2560) : 0
(1552,2240):(4640,2560) : 0
(1374,1884):(1552,2560) : 0
(786,2240):(1374,2560) : 0
(606,1940):(786,2560) : 0
(0,2240):(606,2560) : 0
SEDFFX1
--pins(9)
SI
use :  
dir : i
shape : 
(1462,1066):(1746,1266) : 0
SE
use : �
dir : i
shape : 
(664,1086):(932,1300) : 0
QN
use :  
dir : o
shape : 
(9166,758):(9286,1648) : 0
(9036,758):(9166,866) : 0
(9010,1486):(9166,1648) : 0
(8856,640):(9036,866) : 0
(8854,666):(8856,866) : 0
Q
use : 
dir : o
shape : 
(8600,426):(8722,1784) : 0
(8468,426):(8600,536) : 0
(8590,1674):(8600,1784) : 0
(8468,1674):(8590,1800) : 0
(8168,350):(8468,536) : 0
(8408,1690):(8468,1800) : 0
(8286,1690):(8408,2012) : 0
(8228,1850):(8286,2012) : 0
E
use :  
dir : i
shape : 
(462,1678):(582,1820) : 0
(372,1710):(462,1820) : 0
(250,1710):(372,1962) : 0
(192,1800):(250,1962) : 0
D
use :  
dir : i
shape : 
(2110,1048):(2364,1254) : 0
CK
use : c
dir : i
shape : 
(4900,866):(5148,1084) : 0
VSS
use : g
dir : b
shape : 
(8992,-160):(9400,160) : 0
(8812,-160):(8992,244) : 0
(7908,-160):(8812,160) : 0
(7786,-160):(7908,682) : 0
(6460,-160):(7786,160) : 0
(6280,-160):(6460,436) : 0
(5530,-160):(6280,160) : 0
(5352,-160):(5530,384) : 0
(1714,-160):(5352,160) : 0
(1594,-160):(1714,398) : 0
(348,-160):(1594,160) : 0
(168,-160):(348,244) : 0
(0,-160):(168,160) : 0
VDD
use : p
dir : b
shape : 
(9072,2240):(9400,2560) : 0
(8864,2156):(9072,2560) : 0
(8004,2226):(8864,2560) : 0
(7826,1692):(8004,2560) : 0
(6588,2240):(7826,2560) : 0
(6092,2156):(6588,2560) : 0
(5518,2240):(6092,2560) : 0
(4726,2156):(5518,2560) : 0
(1556,2240):(4726,2560) : 0
(1376,1926):(1556,2560) : 0
(744,2240):(1376,2560) : 0
(564,1972):(744,2560) : 0
(0,2240):(564,2560) : 0
SEDFFHQX4
--pins(8)
SI
use :  
dir : i
shape : 
(742,334):(1024,524) : 0
SE
use : �
dir : i
shape : 
(340,980):(582,1266) : 0
Q
use :  
dir : o
shape : 
(12672,866):(12778,1534) : 0
(12578,690):(12672,1534) : 0
(12492,690):(12578,1466) : 0
E
use : 
dir : i
shape : 
(3548,1098):(3748,1386) : 0
(3408,1110):(3548,1220) : 0
D
use :  
dir : i
shape : 
(2158,866):(2360,1128) : 0
CK
use : c
dir : i
shape : 
(5098,988):(5210,1150) : 0
(4958,988):(5098,1254) : 0
(4842,988):(4958,1150) : 0
VSS
use : g
dir : b
shape : 
(13028,-160):(13200,160) : 0
(12850,-160):(13028,244) : 0
(12292,-160):(12850,160) : 0
(12114,-160):(12292,728) : 0
(11514,-160):(12114,160) : 0
(11334,-160):(11514,244) : 0
(8850,-160):(11334,160) : 0
(8672,-160):(8850,244) : 0
(8050,-160):(8672,160) : 0
(7872,-160):(8050,244) : 0
(6866,-160):(7872,160) : 0
(6686,-160):(6866,574) : 0
(5466,-160):(6686,160) : 0
(5286,-160):(5466,244) : 0
(3644,-160):(5286,160) : 0
(3466,-160):(3644,244) : 0
(2228,-160):(3466,160) : 0
(2050,-160):(2228,244) : 0
(590,-160):(2050,160) : 0
(410,-160):(590,244) : 0
(0,-160):(410,160) : 0
VDD
use : p
dir : b
shape : 
(13034,2240):(13200,2560) : 0
(12856,2156):(13034,2560) : 0
(12292,2240):(12856,2560) : 0
(12114,1470):(12292,2560) : 0
(11514,2240):(12114,2560) : 0
(11060,2156):(11514,2560) : 0
(6440,2240):(11060,2560) : 0
(5956,2156):(6440,2560) : 0
(5402,2240):(5956,2560) : 0
(5224,2156):(5402,2560) : 0
(3636,2240):(5224,2560) : 0
(3458,2156):(3636,2560) : 0
(2224,2240):(3458,2560) : 0
(2044,2156):(2224,2560) : 0
(622,2240):(2044,2560) : 0
(442,2156):(622,2560) : 0
(0,2240):(442,2560) : 0
SEDFFHQX2
--pins(8)
SI
use :  
dir : i
shape : 
(742,334):(1022,524) : 0
SE
use : �
dir : i
shape : 
(340,980):(582,1266) : 0
Q
use : 

dir : o
shape : 
(11724,692):(11726,1466) : 0
(11606,692):(11724,1534) : 0
(11516,692):(11606,854) : 0
(11526,1304):(11606,1534) : 0
(11516,1304):(11526,1466) : 0
E
use : 
dir : i
shape : 
(3544,1098):(3744,1386) : 0
(3404,1110):(3544,1220) : 0
D
use : �
dir : i
shape : 
(2156,866):(2358,1128) : 0
CK
use : c
dir : i
shape : 
(4896,842):(5256,1024) : 0
VSS
use : g
dir : b
shape : 
(11338,-160):(11800,160) : 0
(11158,-160):(11338,244) : 0
(10588,-160):(11158,160) : 0
(10410,-160):(10588,244) : 0
(8800,-160):(10410,160) : 0
(8622,-160):(8800,790) : 0
(8042,-160):(8622,160) : 0
(7864,-160):(8042,684) : 0
(6860,-160):(7864,160) : 0
(6680,-160):(6860,574) : 0
(5460,-160):(6680,160) : 0
(5282,-160):(5460,244) : 0
(3642,-160):(5282,160) : 0
(3462,-160):(3642,244) : 0
(2226,-160):(3462,160) : 0
(2048,-160):(2226,244) : 0
(588,-160):(2048,160) : 0
(410,-160):(588,244) : 0
(0,-160):(410,160) : 0
VDD
use : p
dir : b
shape : 
(11338,2240):(11800,2560) : 0
(11158,2156):(11338,2560) : 0
(10552,2240):(11158,2560) : 0
(10372,2156):(10552,2560) : 0
(6476,2240):(10372,2560) : 0
(6298,2156):(6476,2560) : 0
(5368,2240):(6298,2560) : 0
(5248,1804):(5368,2560) : 0
(3634,2240):(5248,2560) : 0
(3454,2156):(3634,2560) : 0
(2222,2240):(3454,2560) : 0
(2042,2156):(2222,2560) : 0
(620,2240):(2042,2560) : 0
(442,2156):(620,2560) : 0
(0,2240):(442,2560) : 0
SEDFFHQX1
--pins(8)
SI
use :  
dir : i
shape : 
(744,334):(1026,524) : 0
SE
use : �
dir : i
shape : 
(340,980):(584,1266) : 0
Q
use :  
dir : o
shape : 
(10566,648):(10686,1542) : 0
(10454,648):(10566,810) : 0
(10502,1380):(10566,1542) : 0
E
use : 

dir : i
shape : 
(3558,1098):(3758,1386) : 0
(3418,1110):(3558,1220) : 0
D
use :  
dir : i
shape : 
(2164,866):(2368,1128) : 0
CK
use : c
dir : i
shape : 
(4914,842):(5276,1024) : 0
VSS
use : g
dir : b
shape : 
(10338,-160):(10800,160) : 0
(10158,-160):(10338,244) : 0
(9634,-160):(10158,160) : 0
(9454,-160):(9634,244) : 0
(8074,-160):(9454,160) : 0
(7894,-160):(8074,740) : 0
(6844,-160):(7894,160) : 0
(6664,-160):(6844,574) : 0
(5482,-160):(6664,160) : 0
(5302,-160):(5482,244) : 0
(3656,-160):(5302,160) : 0
(3476,-160):(3656,244) : 0
(2236,-160):(3476,160) : 0
(2056,-160):(2236,244) : 0
(592,-160):(2056,160) : 0
(412,-160):(592,244) : 0
(0,-160):(412,160) : 0
VDD
use : p
dir : b
shape : 
(10388,2240):(10800,2560) : 0
(10162,2156):(10388,2560) : 0
(9612,2240):(10162,2560) : 0
(9432,2156):(9612,2560) : 0
(6500,2240):(9432,2560) : 0
(6322,2156):(6500,2560) : 0
(5390,2240):(6322,2560) : 0
(5268,1804):(5390,2560) : 0
(3648,2240):(5268,2560) : 0
(3468,2156):(3648,2560) : 0
(2230,2240):(3468,2560) : 0
(2050,2156):(2230,2560) : 0
(622,2240):(2050,2560) : 0
(444,2156):(622,2560) : 0
(0,2240):(444,2560) : 0
SDFFSHQXL
--pins(8)
SN
use :  
dir : i
shape : 
(7236,1042):(7396,1204) : 0
(7214,1042):(7236,1254) : 0
(7156,1058):(7214,1254) : 0
(7034,1058):(7156,1988) : 0
(4272,1878):(7034,1988) : 0
(4150,1266):(4272,1988) : 0
(4086,1266):(4150,1402) : 0
(3964,1146):(4086,1402) : 0
(3608,1216):(3964,1402) : 0
SI
use : �
dir : i
shape : 
(1514,870):(1728,1070) : 0
(1376,960):(1514,1070) : 0
SE
use :  
dir : i
shape : 
(1764,1180):(1886,1562) : 0
(1636,1400):(1764,1562) : 0
(1286,1452):(1636,1562) : 0
(1232,1412):(1286,1562) : 0
(1110,1228):(1232,1562) : 0
(816,1228):(1110,1338) : 0
(694,1158):(816,1338) : 0
Q
use : 

dir : o
shape : 
(8164,534):(8286,1430) : 0
(8026,534):(8164,696) : 0
(8124,1254):(8164,1430) : 0
(7670,1322):(8124,1430) : 0
(7548,1322):(7670,1648) : 0
(7490,1486):(7548,1648) : 0
D
use :  
dir : i
shape : 
(2336,702):(2344,930) : 0
(2214,702):(2336,988) : 0
(2108,702):(2214,970) : 0
(2062,702):(2108,930) : 0
CK
use : c
dir : i
shape : 
(274,422):(278,584) : 0
(68,324):(274,584) : 0
VSS
use : g
dir : b
shape : 
(7528,-160):(8400,160) : 0
(7348,-160):(7528,650) : 0
(6624,-160):(7348,160) : 0
(6444,-160):(6624,244) : 0
(5040,-160):(6444,160) : 0
(4918,-160):(5040,682) : 0
(3542,-160):(4918,160) : 0
(3362,-160):(3542,372) : 0
(1686,-160):(3362,160) : 0
(1506,-160):(1686,244) : 0
(594,-160):(1506,160) : 0
(414,-160):(594,244) : 0
(0,-160):(414,160) : 0
VDD
use : p
dir : b
shape : 
(8052,2240):(8400,2560) : 0
(7872,1610):(8052,2560) : 0
(7348,2240):(7872,2560) : 0
(7168,2156):(7348,2560) : 0
(6616,2240):(7168,2560) : 0
(6436,2156):(6616,2560) : 0
(4932,2240):(6436,2560) : 0
(4738,2156):(4932,2560) : 0
(4026,2240):(4738,2560) : 0
(3526,2002):(4026,2560) : 0
(1804,2240):(3526,2560) : 0
(1622,2156):(1804,2560) : 0
(584,2240):(1622,2560) : 0
(404,2156):(584,2560) : 0
(0,2240):(404,2560) : 0
SDFFSHQX4
--pins(8)
SN
use :  
dir : i
shape : 
(10264,1072):(10384,1180) : 0
(10086,1072):(10264,1222) : 0
(9384,1112):(10086,1222) : 0
(9360,1074):(9384,1222) : 0
(9238,1074):(9360,2016) : 0
(9164,1074):(9238,1184) : 0
(9174,1788):(9238,2016) : 0
(6726,1908):(9174,2016) : 0
(6604,1680):(6726,2016) : 0
(4394,1680):(6604,1790) : 0
(4394,1412):(4436,1522) : 0
(4272,1380):(4394,1790) : 0
(3750,1380):(4272,1490) : 0
SI
use : �
dir : i
shape : 
(1636,1190):(1674,1352) : 0
(1514,642):(1636,1352) : 0
(1442,642):(1514,752) : 0
(1492,1190):(1514,1352) : 0
SE
use :  
dir : i
shape : 
(912,1146):(936,1292) : 0
(668,1134):(912,1338) : 0
Q
use :  
dir : o
shape : 
(11094,380):(11104,612) : 0
(10972,380):(11094,1516) : 0
(10924,380):(10972,712) : 0
(10776,1408):(10972,1516) : 0
(9746,602):(10924,712) : 0
(10574,1400):(10776,2066) : 0
(10458,1422):(10574,1920) : 0
(10386,1422):(10458,1534) : 0
(9914,1422):(10386,1530) : 0
(9832,1422):(9914,1534) : 0
(9652,1422):(9832,1870) : 0
(9622,502):(9746,712) : 0
(9566,502):(9622,664) : 0
D
use :  
dir : i
shape : 
(2154,658):(2376,1000) : 0
CK
use : c
dir : i
shape : 
(490,836):(662,1020) : 0
(368,836):(490,1110) : 0
VSS
use : g
dir : b
shape : 
(10426,-160):(11200,160) : 0
(10246,-160):(10426,424) : 0
(8346,-160):(10246,160) : 0
(8166,-160):(8346,244) : 0
(6078,-160):(8166,160) : 0
(5896,-160):(6078,580) : 0
(5310,-160):(5896,160) : 0
(5130,-160):(5310,634) : 0
(3566,-160):(5130,160) : 0
(3386,-160):(3566,466) : 0
(1824,-160):(3386,160) : 0
(1644,-160):(1824,244) : 0
(686,-160):(1644,160) : 0
(506,-160):(686,244) : 0
(0,-160):(506,160) : 0
VDD
use : p
dir : b
shape : 
(11060,2240):(11200,2560) : 0
(10938,1688):(11060,2560) : 0
(10234,2240):(10938,2560) : 0
(10054,1688):(10234,2560) : 0
(9408,2240):(10054,2560) : 0
(9228,2156):(9408,2560) : 0
(8628,2240):(9228,2560) : 0
(8448,2156):(8628,2560) : 0
(6146,2240):(8448,2560) : 0
(5966,2156):(6146,2560) : 0
(5338,2240):(5966,2560) : 0
(5158,2156):(5338,2560) : 0
(4560,2240):(5158,2560) : 0
(4380,2156):(4560,2560) : 0
(3754,2240):(4380,2560) : 0
(3574,2156):(3754,2560) : 0
(2018,2240):(3574,2560) : 0
(1838,2008):(2018,2560) : 0
(690,2240):(1838,2560) : 0
(510,2156):(690,2560) : 0
(0,2240):(510,2560) : 0
SDFFSHQX2
--pins(8)
SN
use :  
dir : i
shape : 
(9304,1004):(9426,1788) : 0
(8142,1678):(9304,1788) : 0
(8142,1036):(8178,1198) : 0
(8020,1036):(8142,1788) : 0
(7996,1036):(8020,1198) : 0
(7982,1678):(8020,1788) : 0
(7860,1678):(7982,2050) : 0
(5834,1940):(7860,2050) : 0
(5712,1740):(5834,2050) : 0
(5674,1740):(5712,1946) : 0
(5176,1740):(5674,1850) : 0
(5074,1740):(5176,1946) : 0
(4954,1740):(5074,2078) : 0
(4128,1970):(4954,2078) : 0
(4086,1170):(4128,2078) : 0
(4006,1146):(4086,2078) : 0
(3582,1146):(4006,1278) : 0
(3432,1146):(3582,1324) : 0
(3402,1162):(3432,1324) : 0
SI
use : �
dir : i
shape : 
(1386,1096):(1662,1314) : 0
SE
use : �
dir : i
shape : 
(692,970):(854,1130) : 0
(674,888):(692,1130) : 0
(586,888):(674,1104) : 0
(570,878):(586,1104) : 0
(464,878):(570,998) : 0
Q
use :  
dir : o
shape : 
(9044,614):(9166,1466) : 0
(8986,614):(9044,734) : 0
(8864,1358):(9044,1466) : 0
(8936,614):(8986,724) : 0
(8756,562):(8936,724) : 0
(8686,1358):(8864,1520) : 0
(8514,1358):(8686,1522) : 0
D
use : 
dir : i
shape : 
(1890,870):(2114,1114) : 0
(1864,878):(1890,988) : 0
CK
use : c
dir : i
shape : 
(252,1812):(358,2016) : 0
(114,1812):(252,2054) : 0
(100,1812):(114,2016) : 0
VSS
use : g
dir : b
shape : 
(9614,-160):(9800,160) : 0
(9434,-160):(9614,690) : 0
(7660,-160):(9434,160) : 0
(7480,-160):(7660,244) : 0
(5794,-160):(7480,160) : 0
(5614,-160):(5794,606) : 0
(5000,-160):(5614,160) : 0
(4878,-160):(5000,622) : 0
(3450,-160):(4878,160) : 0
(3270,-160):(3450,428) : 0
(1666,-160):(3270,160) : 0
(1484,-160):(1666,244) : 0
(572,-160):(1484,160) : 0
(392,-160):(572,244) : 0
(0,-160):(392,160) : 0
VDD
use : p
dir : b
shape : 
(9098,2240):(9800,2560) : 0
(8918,1976):(9098,2560) : 0
(8302,2240):(8918,2560) : 0
(8122,1952):(8302,2560) : 0
(5510,2240):(8122,2560) : 0
(5330,1992):(5510,2560) : 0
(3884,2240):(5330,2560) : 0
(3454,2002):(3884,2560) : 0
(1790,2240):(3454,2560) : 0
(1610,2002):(1790,2560) : 0
(578,2240):(1610,2560) : 0
(398,2156):(578,2560) : 0
(0,2240):(398,2560) : 0
SDFFSHQX1
--pins(8)
SN
use :  
dir : i
shape : 
(7464,878):(7586,1000) : 0
(7396,890):(7464,1000) : 0
(7274,890):(7396,1166) : 0
(7214,1004):(7274,1166) : 0
(7156,1058):(7214,1166) : 0
(7034,1058):(7156,1988) : 0
(4272,1878):(7034,1988) : 0
(4150,1266):(4272,1988) : 0
(4086,1266):(4150,1402) : 0
(3964,1146):(4086,1402) : 0
(3608,1216):(3964,1402) : 0
SI
use : �
dir : i
shape : 
(1620,688):(1636,1322) : 0
(1586,688):(1620,1348) : 0
(1514,662):(1586,1348) : 0
(1474,662):(1514,878) : 0
(1440,1186):(1514,1348) : 0
(1406,662):(1474,824) : 0
SE
use :  
dir : i
shape : 
(748,1078):(992,1338) : 0
Q
use :  
dir : o
shape : 
(8164,408):(8286,1430) : 0
(8124,408):(8164,614) : 0
(8124,1254):(8164,1430) : 0
(8056,408):(8124,580) : 0
(7670,1322):(8124,1430) : 0
(7548,1322):(7670,1638) : 0
(7490,1476):(7548,1638) : 0
D
use :  
dir : i
shape : 
(2062,842):(2344,1072) : 0
CK
use : c
dir : i
shape : 
(546,878):(586,988) : 0
(538,878):(546,1130) : 0
(442,878):(538,1134) : 0
(416,878):(442,1196) : 0
(320,1022):(416,1196) : 0
VSS
use : g
dir : b
shape : 
(7506,-160):(8400,160) : 0
(7326,-160):(7506,244) : 0
(6624,-160):(7326,160) : 0
(6444,-160):(6624,244) : 0
(5040,-160):(6444,160) : 0
(4918,-160):(5040,580) : 0
(3542,-160):(4918,160) : 0
(3362,-160):(3542,372) : 0
(1670,-160):(3362,160) : 0
(1490,-160):(1670,244) : 0
(572,-160):(1490,160) : 0
(392,-160):(572,412) : 0
(0,-160):(392,160) : 0
VDD
use : p
dir : b
shape : 
(8052,2240):(8400,2560) : 0
(7872,1610):(8052,2560) : 0
(7360,2240):(7872,2560) : 0
(7180,2156):(7360,2560) : 0
(6616,2240):(7180,2560) : 0
(6436,2156):(6616,2560) : 0
(4932,2240):(6436,2560) : 0
(4738,2156):(4932,2560) : 0
(4026,2240):(4738,2560) : 0
(3526,2002):(4026,2560) : 0
(1972,2240):(3526,2560) : 0
(1850,2004):(1972,2560) : 0
(584,2240):(1850,2560) : 0
(404,2156):(584,2560) : 0
(0,2240):(404,2560) : 0
SDFFSXL
--pins(9)
SN
use :  
dir : i
shape : 
(6374,1934):(6708,2100) : 0
SI
use : �
dir : i
shape : 
(1670,1004):(1736,1254) : 0
(1614,1004):(1670,1262) : 0
(1458,1024):(1614,1262) : 0
SE
use :  
dir : i
shape : 
(440,864):(848,1000) : 0
QN
use :  
dir : o
shape : 
(7530,412):(7652,1880) : 0
(7278,412):(7530,522) : 0
(7424,1772):(7530,1880) : 0
(7236,1772):(7424,1954) : 0
(7156,324):(7278,522) : 0
(7114,1772):(7236,2054) : 0
(7042,324):(7156,486) : 0
Q
use :  
dir : o
shape : 
(7936,1472):(8092,1634) : 0
(7936,596):(8072,758) : 0
(7890,596):(7936,1634) : 0
(7814,622):(7890,1634) : 0
D
use :  
dir : i
shape : 
(2376,990):(2392,1100) : 0
(2174,866):(2376,1120) : 0
CK
use : c
dir : i
shape : 
(74,1348):(400,1534) : 0
VSS
use : g
dir : b
shape : 
(7726,-160):(8400,160) : 0
(7546,-160):(7726,244) : 0
(6820,-160):(7546,160) : 0
(6640,-160):(6820,244) : 0
(6046,-160):(6640,160) : 0
(5866,-160):(6046,244) : 0
(4776,-160):(5866,160) : 0
(4654,-160):(4776,384) : 0
(3702,-160):(4654,160) : 0
(3522,-160):(3702,444) : 0
(1902,-160):(3522,160) : 0
(1720,-160):(1902,244) : 0
(756,-160):(1720,160) : 0
(576,-160):(756,244) : 0
(0,-160):(576,160) : 0
VDD
use : p
dir : b
shape : 
(7820,2240):(8400,2560) : 0
(7608,2156):(7820,2560) : 0
(6952,2240):(7608,2560) : 0
(6952,1420):(7042,1522) : 0
(6862,1420):(6952,2560) : 0
(6830,1446):(6862,2560) : 0
(6252,2240):(6830,2560) : 0
(6072,2002):(6252,2560) : 0
(4922,2240):(6072,2560) : 0
(4740,2002):(4922,2560) : 0
(4224,2240):(4740,2560) : 0
(4102,2002):(4224,2560) : 0
(3510,2240):(4102,2560) : 0
(3330,2156):(3510,2560) : 0
(1848,2240):(3330,2560) : 0
(1726,1982):(1848,2560) : 0
(572,2240):(1726,2560) : 0
(392,2156):(572,2560) : 0
(0,2240):(392,2560) : 0
SDFFSX4
--pins(9)
SN
use :  
dir : i
shape : 
(3802,1924):(4126,2100) : 0
SI
use : �
dir : i
shape : 
(1512,976):(1724,1254) : 0
SE
use :  
dir : i
shape : 
(774,866):(936,1190) : 0
(748,988):(774,1190) : 0
QN
use :  
dir : o
shape : 
(10076,648):(10086,810) : 0
(10076,1304):(10086,1466) : 0
(9896,600):(10076,1466) : 0
(9874,600):(9896,1266) : 0
Q
use :  
dir : o
shape : 
(11046,866):(11126,1534) : 0
(10924,700):(11046,1534) : 0
(10766,700):(10924,810) : 0
(10584,1304):(10924,1466) : 0
(10584,648):(10766,810) : 0
D
use :  
dir : i
shape : 
(2108,876):(2336,1126) : 0
CK
use : c
dir : i
shape : 
(504,1134):(626,1266) : 0
(382,874):(504,1266) : 0
(324,874):(382,1036) : 0
VSS
use : g
dir : b
shape : 
(11104,-160):(11200,160) : 0
(10924,-160):(11104,422) : 0
(10426,-160):(10924,160) : 0
(10246,-160):(10426,422) : 0
(9726,-160):(10246,160) : 0
(9546,-160):(9726,244) : 0
(9010,-160):(9546,160) : 0
(8830,-160):(9010,494) : 0
(7632,-160):(8830,160) : 0
(7450,-160):(7632,244) : 0
(6576,-160):(7450,160) : 0
(6396,-160):(6576,598) : 0
(5218,-160):(6396,160) : 0
(5038,-160):(5218,598) : 0
(3670,-160):(5038,160) : 0
(3490,-160):(3670,580) : 0
(1804,-160):(3490,160) : 0
(1622,-160):(1804,244) : 0
(626,-160):(1622,160) : 0
(446,-160):(626,244) : 0
(0,-160):(446,160) : 0
VDD
use : p
dir : b
shape : 
(11104,2240):(11200,2560) : 0
(10924,1978):(11104,2560) : 0
(10426,2240):(10924,2560) : 0
(10246,1978):(10426,2560) : 0
(9726,2240):(10246,2560) : 0
(9546,2156):(9726,2560) : 0
(8968,2240):(9546,2560) : 0
(8788,1558):(8968,2560) : 0
(8204,2240):(8788,2560) : 0
(8024,1666):(8204,2560) : 0
(7418,2240):(8024,2560) : 0
(7238,1954):(7418,2560) : 0
(6512,2240):(7238,2560) : 0
(6332,1942):(6512,2560) : 0
(5112,2240):(6332,2560) : 0
(4932,1942):(5112,2560) : 0
(4372,2240):(4932,2560) : 0
(4250,1942):(4372,2560) : 0
(3672,2240):(4250,2560) : 0
(3550,2006):(3672,2560) : 0
(1882,2240):(3550,2560) : 0
(1702,2002):(1882,2560) : 0
(396,2240):(1702,2560) : 0
(130,2154):(396,2560) : 0
(0,2240):(130,2560) : 0
SDFFRHQXL
--pins(8)
SI
use :  
dir : i
shape : 
(1754,1134):(1998,1254) : 0
(1602,976):(1754,1254) : 0
(1574,976):(1602,1138) : 0
SE
use : �
dir : i
shape : 
(760,866):(998,1086) : 0
RN
use : �
dir : i
shape : 
(7974,1412):(7982,1522) : 0
(7552,1386):(7974,1552) : 0
Q
use : (
dir : o
shape : 
(8726,604):(8734,1522) : 0
(8610,604):(8726,1930) : 0
(8154,604):(8610,714) : 0
(8562,1412):(8610,1930) : 0
(8512,1770):(8562,1930) : 0
(8032,334):(8154,714) : 0
(7974,334):(8032,496) : 0
D
use :  
dir : i
shape : 
(2070,834):(2390,1004) : 0
CK
use : c
dir : i
shape : 
(466,1034):(590,1254) : 0
(336,1034):(466,1250) : 0
VSS
use : g
dir : b
shape : 
(8582,-160):(8800,160) : 0
(8400,-160):(8582,466) : 0
(7726,-160):(8400,160) : 0
(7224,-160):(7726,244) : 0
(6616,-160):(7224,160) : 0
(6434,-160):(6616,244) : 0
(5030,-160):(6434,160) : 0
(4848,-160):(5030,522) : 0
(3594,-160):(4848,160) : 0
(4288,726):(4346,828) : 0
(4166,576):(4288,828) : 0
(3594,576):(4166,676) : 0
(3414,-160):(3594,676) : 0
(1736,-160):(3414,160) : 0
(1554,-160):(1736,244) : 0
(602,-160):(1554,160) : 0
(422,-160):(602,244) : 0
(0,-160):(422,160) : 0
VDD
use : p
dir : b
shape : 
(8010,2240):(8800,2560) : 0
(7830,1700):(8010,2560) : 0
(6790,2240):(7830,2560) : 0
(6568,2156):(6790,2560) : 0
(5210,2240):(6568,2560) : 0
(5030,2156):(5210,2560) : 0
(3562,2240):(5030,2560) : 0
(3382,1934):(3562,2560) : 0
(1866,2240):(3382,2560) : 0
(1686,1996):(1866,2560) : 0
(490,2240):(1686,2560) : 0
(310,1856):(490,2560) : 0
(0,2240):(310,2560) : 0
SDFFRHQX4
--pins(8)
SI
use :  
dir : i
shape : 
(1458,1342):(1656,1612) : 0
SE
use : �
dir : i
shape : 
(1962,1124):(2180,1234) : 0
(1842,1124):(1962,1254) : 0
(1658,1124):(1842,1234) : 0
(1538,908):(1658,1234) : 0
(1378,908):(1538,1016) : 0
RN
use :  
dir : i
shape : 
(9058,874):(9574,1000) : 0
(9054,874):(9058,984) : 0
Q
use : 

dir : o
shape : 
(12638,1414):(12666,1862) : 0
(12488,1412):(12638,1862) : 0
(12380,1412):(12488,1534) : 0
(12182,698):(12380,1534) : 0
(12014,698):(12182,808) : 0
(11324,1424):(12182,1534) : 0
(11836,358):(12014,808) : 0
(11258,698):(11836,808) : 0
(11146,1414):(11324,1862) : 0
(11110,358):(11258,808) : 0
(11080,358):(11110,804) : 0
D
use :  
dir : i
shape : 
(2088,1412):(2412,1584) : 0
CK
use : c
dir : i
shape : 
(330,952):(580,1254) : 0
VSS
use : g
dir : b
shape : 
(12392,-160):(12800,160) : 0
(12212,-160):(12392,470) : 0
(11636,-160):(12212,160) : 0
(11458,-160):(11636,470) : 0
(10754,-160):(11458,160) : 0
(10632,-160):(10754,720) : 0
(9846,-160):(10632,160) : 0
(9668,-160):(9846,244) : 0
(9070,-160):(9668,160) : 0
(8892,-160):(9070,536) : 0
(6166,-160):(8892,160) : 0
(5988,-160):(6166,598) : 0
(5412,-160):(5988,160) : 0
(5234,-160):(5412,680) : 0
(4534,-160):(5234,160) : 0
(4534,630):(4562,732) : 0
(4414,-160):(4534,732) : 0
(3788,-160):(4414,160) : 0
(4384,630):(4414,732) : 0
(3608,-160):(3788,432) : 0
(2102,-160):(3608,160) : 0
(1924,-160):(2102,244) : 0
(674,-160):(1924,160) : 0
(496,-160):(674,244) : 0
(0,-160):(496,160) : 0
VDD
use : p
dir : b
shape : 
(11996,2240):(12800,2560) : 0
(11818,1820):(11996,2560) : 0
(10624,2240):(11818,2560) : 0
(10504,1484):(10624,2560) : 0
(9762,2240):(10504,2560) : 0
(9584,2156):(9762,2560) : 0
(8900,2240):(9584,2560) : 0
(8722,1978):(8900,2560) : 0
(6282,2240):(8722,2560) : 0
(6104,2156):(6282,2560) : 0
(5482,2240):(6104,2560) : 0
(5362,1964):(5482,2560) : 0
(4736,2240):(5362,2560) : 0
(4558,2156):(4736,2560) : 0
(3746,2240):(4558,2560) : 0
(3566,2156):(3746,2560) : 0
(692,2240):(3566,2560) : 0
(514,2156):(692,2560) : 0
(0,2240):(514,2560) : 0
SDFFRHQX2
--pins(8)
SI
use :  
dir : i
shape : 
(1730,1134):(1968,1258) : 0
(1552,1096):(1730,1258) : 0
SE
use : �
dir : i
shape : 
(766,830):(982,1086) : 0
RN
use : 
dir : i
shape : 
(8432,1264):(8714,1526) : 0
Q
use :  
dir : o
shape : 
(9874,550):(9996,1458) : 0
(9286,550):(9874,660) : 0
(9634,1348):(9874,1458) : 0
(9454,1348):(9634,1920) : 0
(9282,450):(9286,660) : 0
(9102,302):(9282,688) : 0
D
use : �
dir : i
shape : 
(2038,836):(2354,1020) : 0
CK
use : c
dir : i
shape : 
(580,1012):(620,1234) : 0
(460,1012):(580,1254) : 0
(316,1012):(460,1234) : 0
VSS
use : g
dir : b
shape : 
(9680,-160):(10400,160) : 0
(9502,-160):(9680,244) : 0
(8764,-160):(9502,160) : 0
(8270,-160):(8764,244) : 0
(7564,-160):(8270,160) : 0
(7386,-160):(7564,244) : 0
(5508,-160):(7386,160) : 0
(5328,-160):(5508,584) : 0
(3462,-160):(5328,160) : 0
(3340,-160):(3462,656) : 0
(3282,-160):(3340,654) : 0
(1652,-160):(3282,160) : 0
(1474,-160):(1652,244) : 0
(568,-160):(1474,160) : 0
(388,-160):(568,244) : 0
(0,-160):(388,160) : 0
VDD
use : p
dir : b
shape : 
(10306,2240):(10400,2560) : 0
(10126,1600):(10306,2560) : 0
(8914,2240):(10126,2560) : 0
(8734,2156):(8914,2560) : 0
(8178,2240):(8734,2560) : 0
(8000,2156):(8178,2560) : 0
(7556,2240):(8000,2560) : 0
(7324,2156):(7556,2560) : 0
(5518,2240):(7324,2560) : 0
(5340,2156):(5518,2560) : 0
(3508,2240):(5340,2560) : 0
(3330,1994):(3508,2560) : 0
(1838,2240):(3330,2560) : 0
(1660,2002):(1838,2560) : 0
(694,2240):(1660,2560) : 0
(672,2026):(694,2560) : 0
(494,1944):(672,2560) : 0
(472,2026):(494,2560) : 0
(0,2240):(472,2560) : 0
SDFFRHQX1
--pins(8)
SI
use :  
dir : i
shape : 
(1754,1134):(1998,1254) : 0
(1602,976):(1754,1254) : 0
(1574,976):(1602,1138) : 0
SE
use : �
dir : i
shape : 
(760,696):(984,1086) : 0
RN
use : �
dir : i
shape : 
(7600,1386):(8022,1552) : 0
Q
use : �
dir : o
shape : 
(8710,592):(8712,1522) : 0
(8678,592):(8710,1946) : 0
(8590,592):(8678,2042) : 0
(8112,592):(8590,702) : 0
(8562,1412):(8590,2042) : 0
(8496,1658):(8562,2042) : 0
(7990,348):(8112,702) : 0
(7930,348):(7990,510) : 0
D
use :  
dir : i
shape : 
(2070,834):(2390,1004) : 0
CK
use : c
dir : i
shape : 
(336,1034):(590,1254) : 0
VSS
use : g
dir : b
shape : 
(8496,-160):(8800,160) : 0
(8314,-160):(8496,422) : 0
(7704,-160):(8314,160) : 0
(7202,-160):(7704,244) : 0
(6594,-160):(7202,160) : 0
(6414,-160):(6594,244) : 0
(5032,-160):(6414,160) : 0
(4850,-160):(5032,508) : 0
(3552,-160):(4850,160) : 0
(3370,-160):(3552,654) : 0
(1674,-160):(3370,160) : 0
(1494,-160):(1674,244) : 0
(576,-160):(1494,160) : 0
(394,-160):(576,244) : 0
(0,-160):(394,160) : 0
VDD
use : p
dir : b
shape : 
(7994,2240):(8800,2560) : 0
(7814,1714):(7994,2560) : 0
(6790,2240):(7814,2560) : 0
(6568,2156):(6790,2560) : 0
(5256,2240):(6568,2560) : 0
(5034,2156):(5256,2560) : 0
(3562,2240):(5034,2560) : 0
(3382,1926):(3562,2560) : 0
(1866,2240):(3382,2560) : 0
(1686,2002):(1866,2560) : 0
(490,2240):(1686,2560) : 0
(310,1864):(490,2560) : 0
(0,2240):(310,2560) : 0
SDFFRXL
--pins(9)
SI
use :  
dir : i
shape : 
(1948,1104):(2010,1274) : 0
(1768,1104):(1948,1392) : 0
SE
use : �
dir : i
shape : 
(650,858):(960,1090) : 0
RN
use :  
dir : i
shape : 
(3856,1380):(4036,1542) : 0
(3776,1380):(3856,1534) : 0
(3736,1124):(3776,1534) : 0
(3654,1124):(3736,1516) : 0
(3584,1124):(3654,1276) : 0
QN
use :  
dir : o
shape : 
(8890,412):(9012,1922) : 0
(8702,412):(8890,522) : 0
(8810,1666):(8890,1922) : 0
(8744,1812):(8810,1922) : 0
(8564,1812):(8744,2014) : 0
(8522,302):(8702,522) : 0
Q
use :  
dir : o
shape : 
(9618,1724):(9662,1886) : 0
(9496,900):(9618,1886) : 0
(9450,900):(9496,1010) : 0
(9482,1724):(9496,1886) : 0
(9174,566):(9450,1010) : 0
D
use :  
dir : i
shape : 
(2176,750):(2384,1002) : 0
(2140,816):(2176,990) : 0
(2110,828):(2140,990) : 0
CK
use : c
dir : i
shape : 
(334,1292):(626,1534) : 0
VSS
use : g
dir : b
shape : 
(9090,-160):(9800,160) : 0
(8910,-160):(9090,244) : 0
(8236,-160):(8910,160) : 0
(8056,-160):(8236,422) : 0
(7302,-160):(8056,160) : 0
(7122,-160):(7302,498) : 0
(4776,-160):(7122,160) : 0
(5586,604):(5768,808) : 0
(4932,604):(5586,704) : 0
(4776,604):(4932,722) : 0
(4654,-160):(4776,722) : 0
(3706,-160):(4654,160) : 0
(3526,-160):(3706,428) : 0
(1750,-160):(3526,160) : 0
(1570,-160):(1750,244) : 0
(642,-160):(1570,160) : 0
(462,-160):(642,244) : 0
(0,-160):(462,160) : 0
VDD
use : p
dir : b
shape : 
(9254,2240):(9800,2560) : 0
(9074,2156):(9254,2560) : 0
(8342,2240):(9074,2560) : 0
(8162,1978):(8342,2560) : 0
(7268,2240):(8162,2560) : 0
(7088,1972):(7268,2560) : 0
(6030,2240):(7088,2560) : 0
(5532,1972):(6030,2560) : 0
(3908,2240):(5532,2560) : 0
(3728,2156):(3908,2560) : 0
(1978,2240):(3728,2560) : 0
(1798,1972):(1978,2560) : 0
(404,2240):(1798,2560) : 0
(222,2156):(404,2560) : 0
(0,2240):(222,2560) : 0
SDFFRX4
--pins(9)
SI
use :  
dir : i
shape : 
(1492,976):(1672,1326) : 0
(1468,980):(1492,1326) : 0
SE
use : 
dir : i
shape : 
(932,614):(940,1114) : 0
(776,612):(932,1114) : 0
(756,612):(776,1096) : 0
RN
use : #
dir : i
shape : 
(3866,1308):(4108,1664) : 0
QN
use : %
dir : o
shape : 
(10880,570):(11080,1534) : 0
(10870,570):(10880,730) : 0
(10870,1324):(10880,1486) : 0
Q
use :  
dir : o
shape : 
(11724,600):(11778,1486) : 0
(11576,570):(11724,1486) : 0
(11574,570):(11576,988) : 0
(11546,1324):(11576,1486) : 0
(11546,570):(11574,730) : 0
D
use :  
dir : i
shape : 
(2084,1124):(2204,1286) : 0
(2014,1124):(2084,1234) : 0
(1894,878):(2014,1234) : 0
(1856,878):(1894,988) : 0
CK
use : c
dir : i
shape : 
(348,1120):(592,1350) : 0
VSS
use : g
dir : b
shape : 
(12062,-160):(12200,160) : 0
(11884,-160):(12062,422) : 0
(11386,-160):(11884,160) : 0
(11208,-160):(11386,422) : 0
(10710,-160):(11208,160) : 0
(10532,-160):(10710,422) : 0
(9988,-160):(10532,160) : 0
(9808,-160):(9988,422) : 0
(9226,-160):(9808,160) : 0
(9048,-160):(9226,422) : 0
(8456,-160):(9048,160) : 0
(8276,-160):(8456,422) : 0
(7520,-160):(8276,160) : 0
(7342,-160):(7520,484) : 0
(6150,-160):(7342,160) : 0
(6028,-160):(6150,672) : 0
(5170,-160):(6028,160) : 0
(4990,-160):(5170,428) : 0
(4108,-160):(4990,160) : 0
(3930,-160):(4108,606) : 0
(1712,-160):(3930,160) : 0
(1532,-160):(1712,244) : 0
(570,-160):(1532,160) : 0
(390,-160):(570,244) : 0
(0,-160):(390,160) : 0
VDD
use : p
dir : b
shape : 
(12062,2240):(12200,2560) : 0
(11884,1954):(12062,2560) : 0
(11386,2240):(11884,2560) : 0
(11208,1954):(11386,2560) : 0
(10710,2240):(11208,2560) : 0
(10532,1972):(10710,2560) : 0
(9882,2240):(10532,2560) : 0
(9702,1484):(9882,2560) : 0
(8508,2240):(9702,2560) : 0
(8328,1972):(8508,2560) : 0
(7198,2240):(8328,2560) : 0
(7018,1780):(7198,2560) : 0
(5694,2240):(7018,2560) : 0
(5514,1896):(5694,2560) : 0
(3760,2240):(5514,2560) : 0
(3580,2156):(3760,2560) : 0
(2050,2240):(3580,2560) : 0
(1870,1972):(2050,2560) : 0
(448,2240):(1870,2560) : 0
(270,2156):(448,2560) : 0
(0,2240):(270,2560) : 0
SDFFNRX1
--pins(9)
SI
use :  
dir : i
shape : 
(1772,1120):(2016,1362) : 0
SE
use : 
dir : i
shape : 
(648,838):(954,1058) : 0
RN
use : �
dir : i
shape : 
(3780,1590):(4112,1700) : 0
(3658,1138):(3780,1700) : 0
(3572,1138):(3658,1262) : 0
QN
use : "
dir : o
shape : 
(8978,410):(8994,1570) : 0
(8872,410):(8978,1800) : 0
(8778,410):(8872,612) : 0
(8818,1460):(8872,1800) : 0
(8640,1678):(8818,1800) : 0
(8408,410):(8778,520) : 0
(8520,1678):(8640,1900) : 0
(8440,1738):(8520,1900) : 0
Q
use : �
dir : o
shape : 
(9306,604):(9312,1742) : 0
(9176,604):(9306,1874) : 0
(9166,604):(9176,878) : 0
(9126,1488):(9176,1874) : 0
(9126,646):(9166,878) : 0
D
use :  
dir : i
shape : 
(2120,762):(2332,1010) : 0
(2078,770):(2120,1010) : 0
CKN
use : c
dir : i
shape : 
(332,1272):(622,1538) : 0
VSS
use : g
dir : b
shape : 
(9262,-160):(9400,160) : 0
(9084,-160):(9262,244) : 0
(7854,-160):(9084,160) : 0
(7676,-160):(7854,244) : 0
(7052,-160):(7676,160) : 0
(6874,-160):(7052,244) : 0
(4750,-160):(6874,160) : 0
(5686,716):(5744,818) : 0
(5566,604):(5686,818) : 0
(4906,604):(5566,704) : 0
(4750,604):(4906,704) : 0
(4628,-160):(4750,704) : 0
(3688,-160):(4628,160) : 0
(3508,-160):(3688,428) : 0
(1688,-160):(3508,160) : 0
(1508,-160):(1688,244) : 0
(284,-160):(1508,160) : 0
(106,-160):(284,244) : 0
(0,-160):(106,160) : 0
VDD
use : p
dir : b
shape : 
(9258,2240):(9400,2560) : 0
(9026,2156):(9258,2560) : 0
(8240,2240):(9026,2560) : 0
(8060,1754):(8240,2560) : 0
(7196,2240):(8060,2560) : 0
(7016,1968):(7196,2560) : 0
(5998,2240):(7016,2560) : 0
(5502,1968):(5998,2560) : 0
(3850,2240):(5502,2560) : 0
(3672,2156):(3850,2560) : 0
(1968,2240):(3672,2560) : 0
(1788,1972):(1968,2560) : 0
(596,2240):(1788,2560) : 0
(416,2156):(596,2560) : 0
(0,2240):(416,2560) : 0
SDFFNXL
--pins(8)
SI
use :  
dir : i
shape : 
(1438,866):(1688,1000) : 0
(1262,824):(1438,1000) : 0
(1234,824):(1262,934) : 0
SE
use : 
dir : i
shape : 
(1956,1238):(2138,1400) : 0
(1698,1264):(1956,1374) : 0
(1576,1134):(1698,1374) : 0
(1132,1134):(1576,1266) : 0
(1062,1146):(1132,1254) : 0
QN
use :  
dir : o
shape : 
(6940,1674):(7122,1836) : 0
(6932,584):(6952,746) : 0
(6932,1674):(6940,1788) : 0
(6810,584):(6932,1784) : 0
(6770,584):(6810,746) : 0
Q
use :  
dir : o
shape : 
(6274,300):(6454,498) : 0
(6254,974):(6356,1638) : 0
(6220,388):(6274,498) : 0
(6234,974):(6254,1690) : 0
(6220,974):(6234,1084) : 0
(6074,1528):(6234,1690) : 0
(6098,388):(6220,1084) : 0
(5752,612):(6098,722) : 0
D
use :  
dir : i
shape : 
(2266,878):(2352,988) : 0
(2114,670):(2266,988) : 0
(2084,670):(2114,830) : 0
CKN
use : c
dir : i
shape : 
(468,1074):(630,1266) : 0
(428,1048):(468,1266) : 0
(344,1048):(428,1264) : 0
VSS
use : g
dir : b
shape : 
(6896,-160):(7400,160) : 0
(6714,-160):(6896,244) : 0
(6050,-160):(6714,160) : 0
(5868,-160):(6050,244) : 0
(4746,-160):(5868,160) : 0
(4564,-160):(4746,690) : 0
(3490,-160):(4564,160) : 0
(3366,-160):(3490,518) : 0
(1640,-160):(3366,160) : 0
(1458,-160):(1640,244) : 0
(608,-160):(1458,160) : 0
(608,644):(704,746) : 0
(524,-160):(608,746) : 0
(486,-160):(524,720) : 0
(0,-160):(486,160) : 0
VDD
use : p
dir : b
shape : 
(6682,2240):(7400,2560) : 0
(6500,2130):(6682,2560) : 0
(5828,2240):(6500,2560) : 0
(5646,2156):(5828,2560) : 0
(4386,2240):(5646,2560) : 0
(3702,2156):(4386,2560) : 0
(2138,2240):(3702,2560) : 0
(1956,2130):(2138,2560) : 0
(502,2240):(1956,2560) : 0
(282,2156):(502,2560) : 0
(0,2240):(282,2560) : 0
SDFFNX1
--pins(8)
SI
use :  
dir : i
shape : 
(1524,878):(1756,1134) : 0
SE
use : 
dir : i
shape : 
(2108,1324):(2138,1486) : 0
(1956,1252):(2108,1486) : 0
(1334,1252):(1956,1362) : 0
(1180,1134):(1334,1362) : 0
(1132,1134):(1180,1266) : 0
QN
use :  
dir : o
shape : 
(7122,566):(7304,1848) : 0
(7068,1686):(7122,1848) : 0
Q
use :  
dir : o
shape : 
(6810,412):(6932,1628) : 0
(6770,412):(6810,612) : 0
(6338,1520):(6810,1628) : 0
(6556,412):(6770,522) : 0
(6374,346):(6556,522) : 0
(6156,1520):(6338,1680) : 0
D
use :  
dir : i
shape : 
(2280,878):(2352,988) : 0
(2144,670):(2280,988) : 0
(2098,670):(2144,830) : 0
CKN
use : c
dir : i
shape : 
(468,1050):(630,1266) : 0
(344,1024):(468,1266) : 0
VSS
use : g
dir : b
shape : 
(6994,-160):(7400,160) : 0
(6812,-160):(6994,244) : 0
(6150,-160):(6812,160) : 0
(5970,-160):(6150,244) : 0
(4848,-160):(5970,160) : 0
(4666,-160):(4848,718) : 0
(3582,-160):(4666,160) : 0
(3402,-160):(3582,518) : 0
(1704,-160):(3402,160) : 0
(1522,-160):(1704,244) : 0
(672,-160):(1522,160) : 0
(672,670):(816,772) : 0
(550,-160):(672,772) : 0
(0,-160):(550,160) : 0
VDD
use : p
dir : b
shape : 
(6844,2240):(7400,2560) : 0
(6664,2130):(6844,2560) : 0
(5932,2240):(6664,2560) : 0
(5750,2156):(5932,2560) : 0
(4504,2240):(5750,2560) : 0
(4322,2156):(4504,2560) : 0
(2154,2240):(4322,2560) : 0
(1972,2130):(2154,2560) : 0
(392,2240):(1972,2560) : 0
(210,2130):(392,2560) : 0
(0,2240):(210,2560) : 0
SDFFHQXL
--pins(7)
SI
use :  
dir : i
shape : 
(1514,878):(1744,1138) : 0
SE
use : 
dir : i
shape : 
(1920,1252):(2100,1434) : 0
(1326,1252):(1920,1362) : 0
(1172,1134):(1326,1362) : 0
(1124,1134):(1172,1266) : 0
Q
use :  
dir : o
shape : 
(6886,378):(6934,1678) : 0
(6812,378):(6886,1788) : 0
(6764,378):(6812,488) : 0
(6764,1520):(6812,1788) : 0
(6666,334):(6764,488) : 0
(6220,1520):(6764,1680) : 0
(6486,326):(6666,488) : 0
D
use :  
dir : i
shape : 
(2264,878):(2336,988) : 0
(2130,670):(2264,988) : 0
(2084,670):(2130,830) : 0
CK
use : c
dir : i
shape : 
(464,1050):(626,1266) : 0
(342,1024):(464,1266) : 0
VSS
use : g
dir : b
shape : 
(6262,-160):(7000,160) : 0
(6082,-160):(6262,244) : 0
(4748,-160):(6082,160) : 0
(4626,-160):(4748,666) : 0
(3530,-160):(4626,160) : 0
(3408,-160):(3530,518) : 0
(1692,-160):(3408,160) : 0
(1512,-160):(1692,244) : 0
(668,-160):(1512,160) : 0
(668,644):(838,746) : 0
(546,-160):(668,746) : 0
(0,-160):(546,160) : 0
VDD
use : p
dir : b
shape : 
(5976,2240):(7000,2560) : 0
(5796,2156):(5976,2560) : 0
(4474,2240):(5796,2560) : 0
(4292,2156):(4474,2560) : 0
(2302,2240):(4292,2560) : 0
(2122,2130):(2302,2560) : 0
(584,2240):(2122,2560) : 0
(404,2156):(584,2560) : 0
(0,2240):(404,2560) : 0
SDFFHQX4
--pins(7)
SI
use :  
dir : i
shape : 
(1678,866):(1742,1066) : 0
(1500,866):(1678,1092) : 0
(1458,866):(1500,1000) : 0
SE
use : 
dir : i
shape : 
(1852,1186):(2030,1348) : 0
(1380,1202):(1852,1312) : 0
(1258,1134):(1380,1312) : 0
(1054,1134):(1258,1266) : 0
Q
use :  
dir : o
shape : 
(8564,866):(8580,1534) : 0
(8386,650):(8564,1534) : 0
(8382,866):(8386,1534) : 0
(8260,1342):(8382,1504) : 0
D
use :  
dir : i
shape : 
(2300,712):(2312,878) : 0
(2300,1146):(2310,1254) : 0
(2176,712):(2300,1254) : 0
(2134,712):(2176,874) : 0
CK
use : c
dir : i
shape : 
(304,1048):(580,1254) : 0
VSS
use : g
dir : b
shape : 
(8900,-160):(9000,160) : 0
(8722,-160):(8900,430) : 0
(8230,-160):(8722,160) : 0
(8050,-160):(8230,424) : 0
(7442,-160):(8050,160) : 0
(7264,-160):(7442,244) : 0
(6490,-160):(7264,160) : 0
(6370,-160):(6490,574) : 0
(4844,-160):(6370,160) : 0
(4722,-160):(4844,622) : 0
(3534,-160):(4722,160) : 0
(3356,-160):(3534,574) : 0
(1688,-160):(3356,160) : 0
(1510,-160):(1688,244) : 0
(676,-160):(1510,160) : 0
(676,718):(692,820) : 0
(498,-160):(676,820) : 0
(0,-160):(498,160) : 0
VDD
use : p
dir : b
shape : 
(8778,2240):(9000,2560) : 0
(8598,1978):(8778,2560) : 0
(8080,2240):(8598,2560) : 0
(7902,2156):(8080,2560) : 0
(7374,2240):(7902,2560) : 0
(6120,2156):(7374,2560) : 0
(4746,2240):(6120,2560) : 0
(4568,2156):(4746,2560) : 0
(2958,2240):(4568,2560) : 0
(2780,2156):(2958,2560) : 0
(674,2240):(2780,2560) : 0
(496,2156):(674,2560) : 0
(0,2240):(496,2560) : 0
SDFFHQX1
--pins(7)
SI
use :  
dir : i
shape : 
(1474,866):(1848,1096) : 0
SE
use : 
dir : i
shape : 
(1920,1228):(2100,1486) : 0
(1326,1228):(1920,1338) : 0
(1126,1134):(1326,1338) : 0
(1124,1134):(1126,1266) : 0
Q
use :  
dir : o
shape : 
(6886,376):(6934,1678) : 0
(6812,376):(6886,1788) : 0
(6764,376):(6812,486) : 0
(6764,1520):(6812,1788) : 0
(6666,334):(6764,486) : 0
(6200,1520):(6764,1680) : 0
(6486,324):(6666,486) : 0
D
use : 

dir : i
shape : 
(2264,878):(2336,988) : 0
(2130,670):(2264,988) : 0
(2084,670):(2130,830) : 0
CK
use : c
dir : i
shape : 
(464,1050):(626,1266) : 0
(342,1024):(464,1266) : 0
VSS
use : g
dir : b
shape : 
(6262,-160):(7000,160) : 0
(6082,-160):(6262,244) : 0
(4748,-160):(6082,160) : 0
(4626,-160):(4748,666) : 0
(3558,-160):(4626,160) : 0
(3378,-160):(3558,518) : 0
(1692,-160):(3378,160) : 0
(1512,-160):(1692,244) : 0
(668,-160):(1512,160) : 0
(668,644):(812,746) : 0
(546,-160):(668,746) : 0
(0,-160):(546,160) : 0
VDD
use : p
dir : b
shape : 
(6782,2240):(7000,2560) : 0
(6602,2130):(6782,2560) : 0
(5976,2240):(6602,2560) : 0
(5796,2156):(5976,2560) : 0
(4422,2240):(5796,2560) : 0
(3744,2156):(4422,2560) : 0
(2302,2240):(3744,2560) : 0
(2122,2130):(2302,2560) : 0
(584,2240):(2122,2560) : 0
(404,2156):(584,2560) : 0
(0,2240):(404,2560) : 0
SDFFXL
--pins(8)
SI
use :  
dir : i
shape : 
(1430,866):(1676,1000) : 0
(1254,824):(1430,1000) : 0
(1226,824):(1254,934) : 0
SE
use : 
dir : i
shape : 
(1894,1238):(2074,1400) : 0
(1686,1238):(1894,1348) : 0
(1564,1134):(1686,1348) : 0
(1174,1134):(1564,1266) : 0
(994,1116):(1174,1278) : 0
QN
use : 
dir : o
shape : 
(6886,1674):(6904,1836) : 0
(6798,564):(6886,1836) : 0
(6764,520):(6798,1836) : 0
(6618,520):(6764,680) : 0
(6724,1674):(6764,1836) : 0
Q
use :  
dir : o
shape : 
(6350,326):(6354,496) : 0
(6170,300):(6350,496) : 0
(6180,1026):(6278,1638) : 0
(6156,1026):(6180,1690) : 0
(6042,386):(6170,496) : 0
(6042,1026):(6156,1136) : 0
(6000,1528):(6156,1690) : 0
(5920,386):(6042,1136) : 0
(5714,600):(5920,734) : 0
D
use :  
dir : i
shape : 
(2020,628):(2200,988) : 0
(1864,878):(2020,988) : 0
CK
use : c
dir : i
shape : 
(464,1074):(626,1266) : 0
(424,1048):(464,1266) : 0
(342,1048):(424,1264) : 0
VSS
use : g
dir : b
shape : 
(6778,-160):(7000,160) : 0
(6596,-160):(6778,244) : 0
(5948,-160):(6596,160) : 0
(5768,-160):(5948,244) : 0
(4654,-160):(5768,160) : 0
(4474,-160):(4654,690) : 0
(3432,-160):(4474,160) : 0
(3250,-160):(3432,518) : 0
(1628,-160):(3250,160) : 0
(1448,-160):(1628,244) : 0
(604,-160):(1448,160) : 0
(604,644):(700,746) : 0
(520,-160):(604,746) : 0
(482,-160):(520,720) : 0
(0,-160):(482,160) : 0
VDD
use : p
dir : b
shape : 
(6530,2240):(7000,2560) : 0
(6350,2130):(6530,2560) : 0
(5754,2240):(6350,2560) : 0
(5574,2156):(5754,2560) : 0
(4436,2240):(5574,2560) : 0
(3758,2156):(4436,2560) : 0
(2132,2240):(3758,2560) : 0
(1952,2130):(2132,2560) : 0
(584,2240):(1952,2560) : 0
(404,2156):(584,2560) : 0
(0,2240):(404,2560) : 0
OR4X2
--pins(7)
Y
use :  
dir : o
shape : 
(1994,364):(2122,2020) : 0
(1884,364):(1994,750) : 0
(1906,1400):(1994,2020) : 0
D
use : 
dir : i
shape : 
(1456,1400):(1756,1534) : 0
(1328,1104):(1456,1534) : 0
C
use : z
dir : i
shape : 
(812,1054):(1112,1266) : 0
B
use : z
dir : i
shape : 
(444,334):(728,528) : 0
A
use :  
dir : i
shape : 
(78,866):(302,1134) : 0
VSS
use : g
dir : b
shape : 
(1292,-160):(2200,160) : 0
(1102,-160):(1292,244) : 0
(288,-160):(1102,160) : 0
(100,-160):(288,244) : 0
(0,-160):(100,160) : 0
VDD
use : p
dir : b
shape : 
(1672,2240):(2200,2560) : 0
(1484,2156):(1672,2560) : 0
(0,2240):(1484,2560) : 0
OR4X1
--pins(7)
Y
use :  
dir : o
shape : 
(2112,1666):(2122,1842) : 0
(1984,452):(2112,1842) : 0
(1900,452):(1984,614) : 0
(1800,1666):(1984,1842) : 0
D
use : 
dir : i
shape : 
(1508,1110):(1772,1330) : 0
C
use :  
dir : i
shape : 
(972,1110):(1100,1534) : 0
(812,1386):(972,1534) : 0
B
use :  
dir : i
shape : 
(444,1034):(712,1270) : 0
A
use :  
dir : i
shape : 
(78,1312):(312,1546) : 0
VSS
use : g
dir : b
shape : 
(1666,-160):(2200,160) : 0
(1478,-160):(1666,244) : 0
(622,-160):(1478,160) : 0
(434,-160):(622,244) : 0
(0,-160):(434,160) : 0
VDD
use : p
dir : b
shape : 
(1566,2240):(2200,2560) : 0
(1378,2156):(1566,2560) : 0
(0,2240):(1378,2560) : 0
OR3XL
--pins(6)
Y
use :  
dir : o
shape : 
(1582,696):(1708,1742) : 0
(1498,696):(1582,858) : 0
(1516,1412):(1582,1742) : 0
(1430,1580):(1516,1742) : 0
C
use : 
dir : i
shape : 
(796,1274):(1090,1534) : 0
B
use :  
dir : i
shape : 
(436,866):(804,1112) : 0
A
use :  
dir : i
shape : 
(412,1272):(538,2054) : 0
(328,1272):(412,1442) : 0
(118,1946):(412,2054) : 0
VSS
use : g
dir : b
shape : 
(1374,-160):(1800,160) : 0
(1190,-160):(1374,244) : 0
(306,-160):(1190,160) : 0
(120,-160):(306,244) : 0
(0,-160):(120,160) : 0
VDD
use : p
dir : b
shape : 
(1310,2240):(1800,2560) : 0
(1124,2156):(1310,2560) : 0
(0,2240):(1124,2560) : 0
OR3X4
--pins(6)
Y
use :  
dir : o
shape : 
(2414,1358):(2678,1534) : 0
(2414,662):(2548,824) : 0
(2208,662):(2414,1534) : 0
C
use : 
dir : i
shape : 
(1834,826):(1932,936) : 0
(1710,826):(1834,1516) : 0
(1662,1400):(1710,1516) : 0
(1538,1408):(1662,1516) : 0
(1392,1408):(1538,1534) : 0
(1268,1408):(1392,1608) : 0
(472,1498):(1268,1608) : 0
(430,1400):(472,1608) : 0
(308,1208):(430,1608) : 0
(248,1208):(308,1550) : 0
(76,1362):(248,1550) : 0
B
use :  
dir : i
shape : 
(1334,914):(1516,1166) : 0
(596,914):(1334,1024) : 0
(528,878):(596,1024) : 0
(344,862):(528,1024) : 0
A
use :  
dir : i
shape : 
(784,1134):(1096,1388) : 0
VSS
use : g
dir : b
shape : 
(2990,-160):(3200,160) : 0
(2806,-160):(2990,244) : 0
(2098,-160):(2806,160) : 0
(1916,-160):(2098,244) : 0
(1242,-160):(1916,160) : 0
(1058,-160):(1242,444) : 0
(0,-160):(1058,160) : 0
VDD
use : p
dir : b
shape : 
(3020,2240):(3200,2560) : 0
(2836,1966):(3020,2560) : 0
(2306,2240):(2836,2560) : 0
(2122,1966):(2306,2560) : 0
(280,2240):(2122,2560) : 0
(96,2156):(280,2560) : 0
(0,2240):(96,2560) : 0
OR2X4
--pins(5)
Y
use :  
dir : o
shape : 
(1388,648):(1466,810) : 0
(1392,1304):(1400,1466) : 0
(1388,1248):(1392,1466) : 0
(1212,600):(1388,1466) : 0
(1178,600):(1212,1266) : 0
B
use : 
dir : i
shape : 
(686,958):(1022,1326) : 0
A
use :  
dir : i
shape : 
(78,784):(288,1112) : 0
VSS
use : g
dir : b
shape : 
(1844,-160):(2200,160) : 0
(1656,-160):(1844,244) : 0
(1112,-160):(1656,160) : 0
(922,-160):(1112,428) : 0
(288,-160):(922,160) : 0
(100,-160):(288,580) : 0
(0,-160):(100,160) : 0
VDD
use : p
dir : b
shape : 
(1778,2240):(2200,2560) : 0
(1588,2156):(1778,2560) : 0
(1022,2240):(1588,2560) : 0
(834,2156):(1022,2560) : 0
(0,2240):(834,2560) : 0
OR2X2
--pins(5)
Y
use :  
dir : o
shape : 
(1178,392):(1300,1828) : 0
(1096,392):(1178,778) : 0
(1092,1442):(1178,1828) : 0
B
use : 
dir : i
shape : 
(424,828):(674,1116) : 0
A
use :  
dir : i
shape : 
(74,786):(276,1088) : 0
VSS
use : g
dir : b
shape : 
(870,-160):(1400,160) : 0
(690,-160):(870,244) : 0
(276,-160):(690,160) : 0
(96,-160):(276,244) : 0
(0,-160):(96,160) : 0
VDD
use : p
dir : b
shape : 
(870,2240):(1400,2560) : 0
(690,2156):(870,2560) : 0
(0,2240):(690,2560) : 0
OR2X1
--pins(5)
Y
use :  
dir : o
shape : 
(1194,628):(1316,1734) : 0
(1124,628):(1194,790) : 0
(1124,1390):(1194,1734) : 0
(1106,1572):(1124,1734) : 0
B
use : 
dir : i
shape : 
(626,1134):(646,1534) : 0
(456,1134):(626,1542) : 0
(424,1400):(456,1542) : 0
A
use :  
dir : i
shape : 
(84,948):(308,1276) : 0
VSS
use : g
dir : b
shape : 
(738,-160):(1400,160) : 0
(238,-160):(738,244) : 0
(0,-160):(238,160) : 0
VDD
use : p
dir : b
shape : 
(768,2240):(1400,2560) : 0
(580,2118):(768,2560) : 0
(0,2240):(580,2560) : 0
OAI33X1
--pins(9)
Y
use :  
dir : o
shape : 
(2620,1146):(2686,1254) : 0
(2498,536):(2620,1774) : 0
(2386,536):(2498,828) : 0
(1252,1664):(2498,1774) : 0
(1804,720):(2386,828) : 0
(1622,626):(1804,828) : 0
(1072,1638):(1252,1800) : 0
B2
use : 
dir : i
shape : 
(74,928):(282,1266) : 0
B1
use :  
dir : i
shape : 
(464,938):(758,1266) : 0
B0
use :  
dir : i
shape : 
(1082,1074):(1140,1236) : 0
(960,1074):(1082,1522) : 0
(814,1400):(960,1522) : 0
A2
use :  
dir : i
shape : 
(2298,1412):(2336,1522) : 0
(2298,1040):(2328,1202) : 0
(2176,1040):(2298,1522) : 0
(2148,1040):(2176,1202) : 0
A1
use :  
dir : i
shape : 
(1728,1010):(2026,1266) : 0
A0
use :  
dir : i
shape : 
(1564,1412):(1636,1522) : 0
(1442,1072):(1564,1522) : 0
(1344,1072):(1442,1234) : 0
VSS
use : g
dir : b
shape : 
(1040,-160):(2800,160) : 0
(860,-160):(1040,578) : 0
(276,-160):(860,160) : 0
(96,-160):(276,660) : 0
(0,-160):(96,160) : 0
VDD
use : p
dir : b
shape : 
(2434,2240):(2800,2560) : 0
(2254,2156):(2434,2560) : 0
(276,2240):(2254,2560) : 0
(96,1600):(276,2560) : 0
(0,2240):(96,2560) : 0
OAI32X4
--pins(8)
Y
use :  
dir : o
shape : 
(2722,866):(2804,1534) : 0
(2596,696):(2722,1534) : 0
(2422,696):(2596,804) : 0
(2278,1376):(2596,1486) : 0
(2236,642):(2422,804) : 0
(2086,1376):(2278,1538) : 0
B1
use : 
dir : i
shape : 
(76,1134):(284,1480) : 0
B0
use :  
dir : i
shape : 
(436,1910):(782,2098) : 0
A2
use :  
dir : i
shape : 
(1768,1134):(2084,1266) : 0
(1582,1052):(1768,1266) : 0
A1
use :  
dir : i
shape : 
(1390,1412):(1682,1522) : 0
(1266,1054):(1390,1522) : 0
(1206,1054):(1266,1216) : 0
A0
use :  
dir : i
shape : 
(770,1134):(1004,1434) : 0
VSS
use : g
dir : b
shape : 
(2792,-160):(3600,160) : 0
(2608,-160):(2792,244) : 0
(2012,-160):(2608,160) : 0
(1828,-160):(2012,244) : 0
(1396,-160):(1828,160) : 0
(1210,-160):(1396,244) : 0
(0,-160):(1210,160) : 0
VDD
use : p
dir : b
shape : 
(2716,2240):(3600,2560) : 0
(2530,1978):(2716,2560) : 0
(1922,2240):(2530,2560) : 0
(1738,1978):(1922,2560) : 0
(284,2240):(1738,2560) : 0
(98,2156):(284,2560) : 0
(0,2240):(98,2560) : 0
OAI32X1
--pins(8)
Y
use :  
dir : o
shape : 
(2350,720):(2480,1752) : 0
(2308,720):(2350,878) : 0
(1136,1642):(2350,1752) : 0
(1914,720):(2308,828) : 0
(1722,628):(1914,828) : 0
B1
use : 
dir : i
shape : 
(1858,974):(2150,1280) : 0
B0
use :  
dir : i
shape : 
(1598,1412):(1736,1522) : 0
(1468,1084):(1598,1522) : 0
(1406,1084):(1468,1246) : 0
A2
use :  
dir : i
shape : 
(78,1134):(298,1422) : 0
A1
use :  
dir : i
shape : 
(664,912):(804,1022) : 0
(492,912):(664,1254) : 0
A0
use :  
dir : i
shape : 
(864,1226):(1120,1522) : 0
VSS
use : g
dir : b
shape : 
(1104,-160):(2600,160) : 0
(912,-160):(1104,554) : 0
(292,-160):(912,160) : 0
(102,-160):(292,580) : 0
(0,-160):(102,160) : 0
VDD
use : p
dir : b
shape : 
(2070,2240):(2600,2560) : 0
(1880,2130):(2070,2560) : 0
(292,2240):(1880,2560) : 0
(102,2004):(292,2560) : 0
(0,2240):(102,2560) : 0
OAI31X1
--pins(7)
Y
use :  
dir : o
shape : 
(1952,472):(2080,1690) : 0
(1912,472):(1952,612) : 0
(1912,1522):(1952,1690) : 0
(1744,472):(1912,580) : 0
(1144,1580):(1912,1690) : 0
B0
use : 
dir : i
shape : 
(1586,880):(1770,1254) : 0
A2
use :  
dir : i
shape : 
(78,962):(288,1266) : 0
A1
use :  
dir : i
shape : 
(444,866):(822,1014) : 0
A0
use :  
dir : i
shape : 
(972,1098):(1206,1302) : 0
(852,1140):(972,1254) : 0
VSS
use : g
dir : b
shape : 
(1134,-160):(2200,160) : 0
(1112,-160):(1134,174) : 0
(922,-160):(1112,244) : 0
(900,-160):(922,174) : 0
(288,-160):(900,160) : 0
(100,-160):(288,550) : 0
(0,-160):(100,160) : 0
VDD
use : p
dir : b
shape : 
(1644,2240):(2200,2560) : 0
(1456,2156):(1644,2560) : 0
(288,2240):(1456,2560) : 0
(100,1850):(288,2560) : 0
(0,2240):(100,2560) : 0
OAI2BB2X4
--pins(7)
Y
use :  
dir : o
shape : 
(5048,558):(5106,720) : 0
(4926,384):(5048,984) : 0
(2960,384):(4926,492) : 0
(4780,874):(4926,984) : 0
(4580,866):(4780,1652) : 0
(3240,1490):(4580,1652) : 0
(3118,1402):(3240,1652) : 0
(2350,1402):(3118,1512) : 0
(2782,314):(2960,492) : 0
B1
use : 
dir : i
shape : 
(3700,1130):(3816,1240) : 0
(3662,1130):(3700,1258) : 0
(3580,1130):(3662,1292) : 0
(3540,1148):(3580,1292) : 0
(1994,1184):(3540,1292) : 0
(1814,1066):(1994,1292) : 0
B0
use :  
dir : i
shape : 
(4394,912):(4460,1146) : 0
(4272,912):(4394,1254) : 0
(3420,912):(4272,1022) : 0
(3388,912):(3420,1060) : 0
(3296,912):(3388,1074) : 0
(3238,950):(3296,1074) : 0
(2224,964):(3238,1074) : 0
A1N
use :  
dir : i
shape : 
(678,1110):(856,1272) : 0
(578,1110):(678,1266) : 0
(434,1134):(578,1266) : 0
A0N
use :  
dir : i
shape : 
(1342,888):(1492,1050) : 0
(1314,370):(1342,1050) : 0
(1222,370):(1314,998) : 0
(606,370):(1222,478) : 0
(486,370):(606,962) : 0
(460,852):(486,962) : 0
(320,852):(460,1000) : 0
(142,852):(320,1014) : 0
(112,878):(142,988) : 0
VSS
use : g
dir : b
shape : 
(4370,-160):(5200,160) : 0
(4192,-160):(4370,244) : 0
(3654,-160):(4192,160) : 0
(3474,-160):(3654,244) : 0
(2224,-160):(3474,160) : 0
(1462,-160):(2224,244) : 0
(274,-160):(1462,160) : 0
(94,-160):(274,550) : 0
(0,-160):(94,160) : 0
VDD
use : p
dir : b
shape : 
(5084,2240):(5200,2560) : 0
(4906,2156):(5084,2560) : 0
(3990,2240):(4906,2560) : 0
(3810,2156):(3990,2560) : 0
(2896,2240):(3810,2560) : 0
(2718,2156):(2896,2560) : 0
(1836,2240):(2718,2560) : 0
(1658,2156):(1836,2560) : 0
(1046,2240):(1658,2560) : 0
(866,2156):(1046,2560) : 0
(274,2240):(866,2560) : 0
(94,1582):(274,2560) : 0
(0,2240):(94,2560) : 0
OAI2BB2X2
--pins(7)
Y
use :  
dir : o
shape : 
(3358,812):(3482,1846) : 0
(2462,812):(3358,922) : 0
(2632,1736):(3358,1846) : 0
(2446,1736):(2632,1898) : 0
(2338,602):(2462,922) : 0
(1802,1736):(2446,1846) : 0
(2204,602):(2338,712) : 0
(1618,1736):(1802,1898) : 0
B1
use : 
dir : i
shape : 
(3082,1252):(3166,1522) : 0
(3040,1252):(3082,1602) : 0
(2956,1412):(3040,1602) : 0
(2480,1492):(2956,1602) : 0
(2354,1264):(2480,1602) : 0
(2236,1264):(2354,1412) : 0
(1298,1264):(2236,1374) : 0
(1172,1058):(1298,1374) : 0
B0
use :  
dir : i
shape : 
(2740,1274):(2830,1384) : 0
(2616,1040):(2740,1384) : 0
(1840,1040):(2616,1150) : 0
(1716,878):(1840,1150) : 0
(1558,878):(1716,988) : 0
A1N
use :  
dir : i
shape : 
(436,1134):(796,1380) : 0
A0N
use :  
dir : i
shape : 
(76,776):(414,1024) : 0
VSS
use : g
dir : b
shape : 
(3088,-160):(3600,160) : 0
(2902,-160):(3088,244) : 0
(1582,-160):(2902,160) : 0
(1396,-160):(1582,244) : 0
(284,-160):(1396,160) : 0
(98,-160):(284,578) : 0
(0,-160):(98,160) : 0
VDD
use : p
dir : b
shape : 
(3352,2240):(3600,2560) : 0
(3166,2156):(3352,2560) : 0
(2218,2240):(3166,2560) : 0
(2032,2156):(2218,2560) : 0
(1104,2240):(2032,2560) : 0
(920,1804):(1104,2560) : 0
(320,2240):(920,2560) : 0
(134,1664):(320,2560) : 0
(0,2240):(134,2560) : 0
OAI2BB2X1
--pins(7)
Y
use :  
dir : o
shape : 
(2464,878):(2480,988) : 0
(2336,500):(2464,1704) : 0
(2274,500):(2336,662) : 0
(2308,1522):(2336,1704) : 0
(1620,1596):(2308,1704) : 0
B1
use : 
dir : i
shape : 
(1140,1028):(1406,1266) : 0
B0
use : 
dir : i
shape : 
(1536,866):(1778,1190) : 0
A1N
use : �
dir : i
shape : 
(468,1000):(684,1266) : 0
A0N
use :  
dir : i
shape : 
(78,784):(338,1014) : 0
VSS
use : g
dir : b
shape : 
(1654,-160):(2600,160) : 0
(1464,-160):(1654,424) : 0
(292,-160):(1464,160) : 0
(102,-160):(292,244) : 0
(0,-160):(102,160) : 0
VDD
use : p
dir : b
shape : 
(2240,2240):(2600,2560) : 0
(2048,2156):(2240,2560) : 0
(1126,2240):(2048,2560) : 0
(934,2156):(1126,2560) : 0
(394,2240):(934,2560) : 0
(362,2156):(394,2560) : 0
(234,2130):(362,2560) : 0
(202,2156):(234,2560) : 0
(0,2240):(202,2560) : 0
OAI2BB1X4
--pins(6)
Y
use :  
dir : o
shape : 
(3240,340):(3338,502) : 0
(3164,340):(3240,1242) : 0
(3122,340):(3164,1800) : 0
(3114,366):(3122,1800) : 0
(2640,366):(3114,476) : 0
(2956,1134):(3114,1800) : 0
(2278,1402):(2956,1512) : 0
(2618,340):(2640,476) : 0
(2432,340):(2618,502) : 0
(2032,1376):(2278,1538) : 0
(1558,1402):(2032,1512) : 0
(1520,1402):(1558,1538) : 0
(1334,1376):(1520,1538) : 0
B0
use : 
dir : i
shape : 
(1156,1078):(1648,1266) : 0
A1N
use :  
dir : i
shape : 
(76,962):(284,1266) : 0
A0N
use :  
dir : i
shape : 
(662,1078):(1004,1266) : 0
VSS
use : g
dir : b
shape : 
(1680,-160):(3600,160) : 0
(1494,-160):(1680,424) : 0
(982,-160):(1494,160) : 0
(796,-160):(982,424) : 0
(0,-160):(796,160) : 0
VDD
use : p
dir : b
shape : 
(2566,2240):(3600,2560) : 0
(2380,1754):(2566,2560) : 0
(1868,2240):(2380,2560) : 0
(1682,1754):(1868,2560) : 0
(1134,2240):(1682,2560) : 0
(950,1888):(1134,2560) : 0
(284,2240):(950,2560) : 0
(98,1494):(284,2560) : 0
(0,2240):(98,2560) : 0
OAI2BB1X2
--pins(6)
Y
use :  
dir : o
shape : 
(2066,584):(2108,1254) : 0
(1978,584):(2066,1462) : 0
(1778,584):(1978,692) : 0
(1936,1146):(1978,1462) : 0
(1834,1352):(1936,1462) : 0
(1644,1352):(1834,1514) : 0
(1588,530):(1778,692) : 0
B0
use : 
dir : i
shape : 
(1070,758):(1406,1014) : 0
A1N
use :  
dir : i
shape : 
(120,800):(330,1066) : 0
A0N
use :  
dir : i
shape : 
(846,1134):(1136,1266) : 0
(718,1084):(846,1266) : 0
VSS
use : g
dir : b
shape : 
(2498,-160):(2600,160) : 0
(2308,-160):(2498,578) : 0
(1036,-160):(2308,160) : 0
(844,-160):(1036,578) : 0
(0,-160):(844,160) : 0
VDD
use : p
dir : b
shape : 
(2218,2240):(2600,2560) : 0
(2026,2156):(2218,2560) : 0
(1474,2240):(2026,2560) : 0
(1284,1944):(1474,2560) : 0
(596,2240):(1284,2560) : 0
(406,2156):(596,2560) : 0
(0,2240):(406,2560) : 0
OAI2BB1X1
--pins(6)
Y
use :  
dir : o
shape : 
(1596,686):(1720,1826) : 0
(1516,686):(1596,848) : 0
(1558,1678):(1596,1826) : 0
(1356,1716):(1558,1826) : 0
(1170,1716):(1356,1878) : 0
B0
use : 
dir : i
shape : 
(796,1052):(1132,1280) : 0
A1N
use :  
dir : i
shape : 
(284,1224):(370,1386) : 0
(76,1224):(284,1534) : 0
A0N
use :  
dir : i
shape : 
(340,848):(644,1064) : 0
VSS
use : g
dir : b
shape : 
(1026,-160):(1800,160) : 0
(840,-160):(1026,244) : 0
(0,-160):(840,160) : 0
VDD
use : p
dir : b
shape : 
(1660,2240):(1800,2560) : 0
(1630,2156):(1660,2560) : 0
(1506,2130):(1630,2560) : 0
(1476,2156):(1506,2560) : 0
(938,2240):(1476,2560) : 0
(98,2156):(938,2560) : 0
(0,2240):(98,2560) : 0
OAI22X4
--pins(7)
Y
use :  
dir : o
shape : 
(4880,866):(4924,1534) : 0
(4756,316):(4880,1534) : 0
(2652,316):(4756,426) : 0
(4718,866):(4756,1534) : 0
(4458,1404):(4718,1514) : 0
(4274,1404):(4458,1854) : 0
(4170,1404):(4274,1534) : 0
(3074,1404):(4170,1514) : 0
(2890,1404):(3074,1854) : 0
(2740,1404):(2890,1534) : 0
(1688,1404):(2740,1514) : 0
(1504,1404):(1688,1854) : 0
(304,1404):(1504,1514) : 0
(120,1404):(304,1852) : 0
B1
use : 
dir : i
shape : 
(2064,1074):(2188,1278) : 0
(1134,1170):(2064,1278) : 0
(952,1100):(1134,1278) : 0
(830,1100):(952,1254) : 0
(682,1100):(830,1210) : 0
B0
use :  
dir : i
shape : 
(1520,898):(1840,1060) : 0
(1374,880):(1520,1060) : 0
(240,880):(1374,990) : 0
(116,880):(240,1254) : 0
A1
use :  
dir : i
shape : 
(3814,898):(3874,1060) : 0
(3690,880):(3814,1060) : 0
(2706,880):(3690,990) : 0
(2706,1126):(2740,1254) : 0
(2616,880):(2706,1254) : 0
(2582,880):(2616,1236) : 0
(2398,1074):(2582,1236) : 0
A0
use :  
dir : i
shape : 
(4234,1074):(4358,1278) : 0
(4170,1134):(4234,1278) : 0
(3496,1170):(4170,1278) : 0
(3372,1100):(3496,1278) : 0
(3330,1100):(3372,1254) : 0
(2988,1100):(3330,1210) : 0
VSS
use : g
dir : b
shape : 
(2056,-160):(5000,160) : 0
(1872,-160):(2056,422) : 0
(1364,-160):(1872,160) : 0
(1180,-160):(1364,422) : 0
(670,-160):(1180,160) : 0
(488,-160):(670,422) : 0
(0,-160):(488,160) : 0
VDD
use : p
dir : b
shape : 
(3766,2240):(5000,2560) : 0
(3582,1864):(3766,2560) : 0
(2380,2240):(3582,2560) : 0
(2196,1864):(2380,2560) : 0
(996,2240):(2196,2560) : 0
(812,1864):(996,2560) : 0
(0,2240):(812,2560) : 0
OAI22X1
--pins(7)
Y
use :  
dir : o
shape : 
(1952,716):(2080,1788) : 0
(1912,716):(1952,878) : 0
(1022,1678):(1952,1788) : 0
(1534,716):(1912,826) : 0
(1406,626):(1534,826) : 0
(1344,626):(1406,788) : 0
(834,1652):(1022,1814) : 0
B1
use : 
dir : i
shape : 
(78,1134):(466,1310) : 0
B0
use :  
dir : i
shape : 
(700,866):(888,1040) : 0
(444,866):(700,1022) : 0
A1
use :  
dir : i
shape : 
(1544,1170):(1756,1534) : 0
A0
use :  
dir : i
shape : 
(1150,946):(1388,1266) : 0
VSS
use : g
dir : b
shape : 
(712,-160):(2200,160) : 0
(522,-160):(712,244) : 0
(0,-160):(522,160) : 0
VDD
use : p
dir : b
shape : 
(1756,2240):(2200,2560) : 0
(1566,2156):(1756,2560) : 0
(288,2240):(1566,2560) : 0
(100,2156):(288,2560) : 0
(0,2240):(100,2560) : 0
OAI222XL
--pins(9)
Y
use :  
dir : o
shape : 
(2564,838):(2686,1788) : 0
(2376,838):(2564,948) : 0
(2296,1678):(2564,1788) : 0
(2302,722):(2376,948) : 0
(2180,562):(2302,948) : 0
(2116,1658):(2296,1820) : 0
(2122,562):(2180,724) : 0
(1986,1666):(2116,1800) : 0
(870,1684):(1986,1792) : 0
(690,1658):(870,1820) : 0
C1
use : 
dir : i
shape : 
(1720,1014):(2026,1266) : 0
C0
use :  
dir : i
shape : 
(2172,1230):(2428,1534) : 0
B1
use :  
dir : i
shape : 
(74,1134):(276,1430) : 0
B0
use :  
dir : i
shape : 
(424,826):(674,1116) : 0
A1
use :  
dir : i
shape : 
(1124,1154):(1352,1536) : 0
A0
use :  
dir : i
shape : 
(706,1278):(976,1534) : 0
VSS
use : g
dir : b
shape : 
(870,-160):(2800,160) : 0
(690,-160):(870,244) : 0
(276,-160):(690,160) : 0
(96,-160):(276,244) : 0
(0,-160):(96,160) : 0
VDD
use : p
dir : b
shape : 
(1582,2240):(2800,2560) : 0
(1402,2156):(1582,2560) : 0
(276,2240):(1402,2560) : 0
(96,2156):(276,2560) : 0
(0,2240):(96,2560) : 0
OAI221XL
--pins(8)
Y
use :  
dir : o
shape : 
(2350,516):(2480,1840) : 0
(2190,516):(2350,678) : 0
(1980,1730):(2350,1840) : 0
(1790,1730):(1980,1892) : 0
(922,1730):(1790,1840) : 0
(732,1730):(922,1892) : 0
C0
use : 
dir : i
shape : 
(1936,1042):(2150,1308) : 0
B1
use :  
dir : i
shape : 
(78,1280):(292,1642) : 0
B0
use :  
dir : i
shape : 
(374,866):(718,1100) : 0
A1
use :  
dir : i
shape : 
(1606,1400):(1736,1522) : 0
(1436,1400):(1606,1510) : 0
(1244,1278):(1436,1510) : 0
A0
use :  
dir : i
shape : 
(1032,1284):(1038,1558) : 0
(842,1280):(1032,1558) : 0
(672,1284):(842,1558) : 0
VSS
use : g
dir : b
shape : 
(922,-160):(2600,160) : 0
(732,-160):(922,244) : 0
(292,-160):(732,160) : 0
(102,-160):(292,244) : 0
(0,-160):(102,160) : 0
VDD
use : p
dir : b
shape : 
(1554,2240):(2600,2560) : 0
(1362,2156):(1554,2560) : 0
(292,2240):(1362,2560) : 0
(102,2156):(292,2560) : 0
(0,2240):(102,2560) : 0
OAI221X4
--pins(8)
Y
use :  
dir : o
shape : 
(3480,866):(3560,1534) : 0
(3416,580):(3480,1534) : 0
(3364,308):(3416,1534) : 0
(3352,308):(3364,1950) : 0
(3228,308):(3352,692) : 0
(3350,866):(3352,1950) : 0
(3176,1340):(3350,1950) : 0
C0
use : 
dir : i
shape : 
(1896,1120):(2104,1392) : 0
B1
use :  
dir : i
shape : 
(78,1308):(330,1580) : 0
B0
use :  
dir : i
shape : 
(440,814):(810,1034) : 0
A1
use :  
dir : i
shape : 
(1574,1146):(1700,1266) : 0
(1408,1158):(1574,1266) : 0
(1280,1158):(1408,1470) : 0
(1220,1308):(1280,1470) : 0
A0
use :  
dir : i
shape : 
(804,1302):(1036,1578) : 0
VSS
use : g
dir : b
shape : 
(3812,-160):(4000,160) : 0
(3626,-160):(3812,646) : 0
(3020,-160):(3626,160) : 0
(2832,-160):(3020,648) : 0
(904,-160):(2832,160) : 0
(716,-160):(904,244) : 0
(286,-160):(716,160) : 0
(100,-160):(286,244) : 0
(0,-160):(100,160) : 0
VDD
use : p
dir : b
shape : 
(3760,2240):(4000,2560) : 0
(3574,1752):(3760,2560) : 0
(2944,2240):(3574,2560) : 0
(2758,2156):(2944,2560) : 0
(2328,2240):(2758,2560) : 0
(2140,2156):(2328,2560) : 0
(1520,2240):(2140,2560) : 0
(1334,2156):(1520,2560) : 0
(286,2240):(1334,2560) : 0
(100,2156):(286,2560) : 0
(0,2240):(100,2560) : 0
OAI221X2
--pins(8)
Y
use :  
dir : o
shape : 
(3952,690):(4064,1660) : 0
(3940,636):(3952,1660) : 0
(3828,636):(3940,880) : 0
(3464,1550):(3940,1660) : 0
(3432,1550):(3464,1678) : 0
(3308,1550):(3432,1808) : 0
(3248,1646):(3308,1808) : 0
(2338,1678):(3248,1788) : 0
(2156,1678):(2338,1840) : 0
(2006,1678):(2156,1800) : 0
(966,1678):(2006,1788) : 0
(782,1678):(966,1840) : 0
C0
use : 
dir : i
shape : 
(3294,1134):(3806,1266) : 0
B1
use :  
dir : i
shape : 
(408,1104):(1480,1214) : 0
(226,1092):(408,1254) : 0
(116,1146):(226,1254) : 0
B0
use :  
dir : i
shape : 
(946,1324):(1094,1486) : 0
(822,1324):(946,1522) : 0
(654,1324):(822,1486) : 0
A1
use :  
dir : i
shape : 
(2638,1124):(3024,1234) : 0
(2514,1104):(2638,1234) : 0
(2008,1104):(2514,1214) : 0
(1908,1104):(2008,1254) : 0
(1884,1104):(1908,1280) : 0
(1726,1120):(1884,1280) : 0
A0
use :  
dir : i
shape : 
(2392,1400):(2480,1534) : 0
(2208,1324):(2392,1534) : 0
(2048,1400):(2208,1534) : 0
VSS
use : g
dir : b
shape : 
(1738,-160):(4600,160) : 0
(1554,-160):(1738,422) : 0
(966,-160):(1554,160) : 0
(782,-160):(966,422) : 0
(278,-160):(782,160) : 0
(96,-160):(278,422) : 0
(0,-160):(96,160) : 0
VDD
use : p
dir : b
shape : 
(3818,2240):(4600,2560) : 0
(3634,1800):(3818,2560) : 0
(3024,2240):(3634,2560) : 0
(2842,1968):(3024,2560) : 0
(1652,2240):(2842,2560) : 0
(1468,1968):(1652,2560) : 0
(278,2240):(1468,2560) : 0
(96,1858):(278,2560) : 0
(0,2240):(96,2560) : 0
OAI221X1
--pins(8)
Y
use :  
dir : o
shape : 
(2620,1658):(2716,1820) : 0
(2498,564):(2620,1820) : 0
(2408,564):(2498,726) : 0
(796,1658):(2498,1820) : 0
C0
use : 
dir : i
shape : 
(2034,1066):(2376,1280) : 0
B1
use :  
dir : i
shape : 
(74,1134):(446,1310) : 0
B0
use :  
dir : i
shape : 
(424,798):(824,1000) : 0
A1
use :  
dir : i
shape : 
(1346,1134):(1676,1342) : 0
A0
use :  
dir : i
shape : 
(750,1120):(1162,1346) : 0
VSS
use : g
dir : b
shape : 
(1082,-160):(2800,160) : 0
(902,-160):(1082,244) : 0
(276,-160):(902,160) : 0
(96,-160):(276,244) : 0
(0,-160):(96,160) : 0
VDD
use : p
dir : b
shape : 
(1676,2240):(2800,2560) : 0
(1646,2156):(1676,2560) : 0
(1524,2130):(1646,2560) : 0
(1496,2156):(1524,2560) : 0
(276,2240):(1496,2560) : 0
(96,2156):(276,2560) : 0
(0,2240):(96,2560) : 0
OAI21XL
--pins(6)
Y
use :  
dir : o
shape : 
(1286,878):(1300,1830) : 0
(1178,322):(1286,1830) : 0
(1164,322):(1178,988) : 0
(954,1722):(1178,1830) : 0
(1092,322):(1164,430) : 0
(774,1696):(954,1858) : 0
B0
use : 
dir : i
shape : 
(774,1280):(1056,1534) : 0
A1
use :  
dir : i
shape : 
(96,866):(276,1236) : 0
A0
use :  
dir : i
shape : 
(586,958):(776,1142) : 0
(464,878):(586,1142) : 0
(424,958):(464,1142) : 0
VSS
use : g
dir : b
shape : 
(572,-160):(1400,160) : 0
(392,-160):(572,244) : 0
(0,-160):(392,160) : 0
VDD
use : p
dir : b
shape : 
(1252,2240):(1400,2560) : 0
(1072,2156):(1252,2560) : 0
(276,2240):(1072,2560) : 0
(96,1820):(276,2560) : 0
(0,2240):(96,2560) : 0
OAI21X4
--pins(6)
Y
use :  
dir : o
shape : 
(3560,626):(3618,880) : 0
(3430,626):(3560,1534) : 0
(3350,662):(3430,1534) : 0
(2658,662):(3350,772) : 0
(3152,1416):(3350,1526) : 0
(2964,1390):(3152,1552) : 0
(2446,1416):(2964,1526) : 0
(2386,1390):(2446,1552) : 0
(2258,1390):(2386,1730) : 0
(992,1622):(2258,1730) : 0
(804,1596):(992,1758) : 0
B0
use : 
dir : i
shape : 
(2524,1120):(2976,1280) : 0
A1
use :  
dir : i
shape : 
(1576,1100):(1874,1210) : 0
(1504,1100):(1576,1266) : 0
(1378,1100):(1504,1486) : 0
(418,1376):(1378,1486) : 0
(292,1066):(418,1486) : 0
(262,1066):(292,1266) : 0
(232,1066):(262,1254) : 0
(118,1146):(232,1254) : 0
A0
use :  
dir : i
shape : 
(2182,1010):(2242,1172) : 0
(2056,880):(2182,1172) : 0
(1168,880):(2056,990) : 0
(1042,880):(1168,1228) : 0
(984,1066):(1042,1228) : 0
(846,1066):(984,1254) : 0
(672,1066):(846,1228) : 0
VSS
use : g
dir : b
shape : 
(2094,-160):(4000,160) : 0
(1906,-160):(2094,422) : 0
(1388,-160):(1906,160) : 0
(1202,-160):(1388,422) : 0
(684,-160):(1202,160) : 0
(496,-160):(684,422) : 0
(0,-160):(496,160) : 0
VDD
use : p
dir : b
shape : 
(3506,2240):(4000,2560) : 0
(3320,1766):(3506,2560) : 0
(2798,2240):(3320,2560) : 0
(2612,1766):(2798,2560) : 0
(1720,2240):(2612,2560) : 0
(1532,1894):(1720,2560) : 0
(286,2240):(1532,2560) : 0
(100,1694):(286,2560) : 0
(0,2240):(100,2560) : 0
OAI21X2
--pins(6)
Y
use :  
dir : o
shape : 
(2566,622):(2686,1840) : 0
(2564,622):(2566,1892) : 0
(2228,622):(2564,730) : 0
(2302,1730):(2564,1892) : 0
(1676,1730):(2302,1840) : 0
(2106,526):(2228,730) : 0
(2046,526):(2106,688) : 0
(1496,1730):(1676,1892) : 0
(276,1730):(1496,1840) : 0
(96,1730):(276,1892) : 0
B0
use : 
dir : i
shape : 
(1750,1102):(2358,1264) : 0
A1
use :  
dir : i
shape : 
(976,1228):(1124,1390) : 0
(946,1228):(976,1414) : 0
(814,1228):(946,1522) : 0
(646,1228):(814,1414) : 0
A0
use :  
dir : i
shape : 
(1422,1210):(1480,1372) : 0
(1300,920):(1422,1372) : 0
(464,920):(1300,1028) : 0
(238,866):(464,1028) : 0
(236,878):(238,1028) : 0
(114,878):(236,988) : 0
VSS
use : g
dir : b
shape : 
(1464,-160):(2800,160) : 0
(1284,-160):(1464,560) : 0
(678,-160):(1284,160) : 0
(498,-160):(678,244) : 0
(0,-160):(498,160) : 0
VDD
use : p
dir : b
shape : 
(2078,2240):(2800,2560) : 0
(1898,2156):(2078,2560) : 0
(976,2240):(1898,2560) : 0
(796,2156):(976,2560) : 0
(0,2240):(796,2560) : 0
OAI21X1
--pins(6)
Y
use :  
dir : o
shape : 
(1560,588):(1682,1830) : 0
(1558,536):(1560,1830) : 0
(1320,536):(1558,698) : 0
(1026,1722):(1558,1830) : 0
(840,1696):(1026,1858) : 0
B0
use : 
dir : i
shape : 
(1108,1120):(1364,1408) : 0
(1102,1120):(1108,1280) : 0
A1
use :  
dir : i
shape : 
(328,866):(480,1000) : 0
(142,852):(328,1014) : 0
(76,866):(142,1000) : 0
A0
use :  
dir : i
shape : 
(436,1134):(850,1266) : 0
VSS
use : g
dir : b
shape : 
(698,-160):(1800,160) : 0
(512,-160):(698,244) : 0
(0,-160):(512,160) : 0
VDD
use : p
dir : b
shape : 
(1440,2240):(1800,2560) : 0
(1254,2156):(1440,2560) : 0
(284,2240):(1254,2560) : 0
(98,1810):(284,2560) : 0
(0,2240):(98,2560) : 0
OAI211X4
--pins(7)
Y
use :  
dir : o
shape : 
(3104,600):(3124,1266) : 0
(2920,600):(3104,1514) : 0
(2576,636):(2920,798) : 0
(2402,1352):(2920,1514) : 0
C0
use : 
dir : i
shape : 
(738,852):(1120,1014) : 0
B0
use :  
dir : i
shape : 
(1346,1074):(1702,1324) : 0
A1
use :  
dir : i
shape : 
(674,1138):(732,1300) : 0
(550,1138):(674,1522) : 0
(472,1412):(550,1522) : 0
A0
use :  
dir : i
shape : 
(76,1022):(372,1270) : 0
VSS
use : g
dir : b
shape : 
(3104,-160):(3200,160) : 0
(2920,-160):(3104,422) : 0
(2414,-160):(2920,160) : 0
(2230,-160):(2414,422) : 0
(636,-160):(2230,160) : 0
(452,-160):(636,244) : 0
(0,-160):(452,160) : 0
VDD
use : p
dir : b
shape : 
(2930,2240):(3200,2560) : 0
(2748,1944):(2930,2560) : 0
(2242,2240):(2748,2560) : 0
(2058,1944):(2242,2560) : 0
(1400,2240):(2058,2560) : 0
(808,2156):(1400,2560) : 0
(0,2240):(808,2560) : 0
OAI211X2
--pins(7)
Y
use :  
dir : o
shape : 
(3262,620):(3388,1510) : 0
(2638,620):(3262,728) : 0
(3122,1400):(3262,1510) : 0
(3082,1400):(3122,1522) : 0
(2998,1400):(3082,1840) : 0
(2956,1412):(2998,1840) : 0
(2640,1730):(2956,1840) : 0
(2368,1730):(2640,1892) : 0
(2596,612):(2638,728) : 0
(2410,566):(2596,728) : 0
(1724,1730):(2368,1840) : 0
(1538,1730):(1724,1904) : 0
(284,1730):(1538,1840) : 0
(98,1730):(284,1892) : 0
C0
use : 
dir : i
shape : 
(3076,838):(3136,1000) : 0
(2950,838):(3076,1254) : 0
(2026,1146):(2950,1254) : 0
(1900,920):(2026,1254) : 0
B0
use :  
dir : i
shape : 
(2728,878):(2762,988) : 0
(2280,852):(2728,1014) : 0
A1
use :  
dir : i
shape : 
(1004,1228):(1156,1390) : 0
(974,1228):(1004,1414) : 0
(838,1228):(974,1522) : 0
(666,1228):(838,1414) : 0
A0
use :  
dir : i
shape : 
(1462,1210):(1522,1372) : 0
(1336,920):(1462,1372) : 0
(478,920):(1336,1028) : 0
(430,866):(478,1028) : 0
(246,852):(430,1028) : 0
(242,878):(246,1028) : 0
(118,878):(242,988) : 0
VSS
use : g
dir : b
shape : 
(1506,-160):(3600,160) : 0
(1320,-160):(1506,560) : 0
(698,-160):(1320,160) : 0
(512,-160):(698,244) : 0
(0,-160):(512,160) : 0
VDD
use : p
dir : b
shape : 
(2138,2240):(3600,2560) : 0
(1952,2156):(2138,2560) : 0
(1004,2240):(1952,2560) : 0
(818,2156):(1004,2560) : 0
(0,2240):(818,2560) : 0
OAI211X1
--pins(7)
Y
use :  
dir : o
shape : 
(1956,596):(2080,1804) : 0
(1952,542):(1956,1858) : 0
(1678,542):(1952,704) : 0
(1700,1696):(1952,1858) : 0
(1044,1696):(1700,1804) : 0
(856,1696):(1044,1858) : 0
C0
use : 
dir : i
shape : 
(1128,1120):(1388,1408) : 0
(1122,1120):(1128,1280) : 0
B0
use :  
dir : i
shape : 
(1544,866):(1756,1204) : 0
A1
use :  
dir : i
shape : 
(334,866):(488,1000) : 0
(144,852):(334,1014) : 0
(78,866):(144,1000) : 0
A0
use :  
dir : i
shape : 
(444,1134):(866,1266) : 0
VSS
use : g
dir : b
shape : 
(712,-160):(2200,160) : 0
(522,-160):(712,244) : 0
(0,-160):(522,160) : 0
VDD
use : p
dir : b
shape : 
(1466,2240):(2200,2560) : 0
(1278,2156):(1466,2560) : 0
(288,2240):(1278,2560) : 0
(100,1810):(288,2560) : 0
(0,2240):(100,2560) : 0
NOR4BBX1
--pins(7)
Y
use :  
dir : o
shape : 
(2614,384):(2736,1788) : 0
(1776,384):(2614,492) : 0
(2028,1678):(2614,1788) : 0
(1848,1678):(2028,1840) : 0
(1626,384):(1776,678) : 0
(1596,446):(1626,678) : 0
(836,446):(1596,608) : 0
D
use : 
dir : i
shape : 
(806,1146):(936,1254) : 0
(684,786):(806,1254) : 0
C
use : z
dir : i
shape : 
(1240,1146):(1286,1254) : 0
(1118,824):(1240,1254) : 0
(1010,824):(1118,986) : 0
BN
use :  
dir : i
shape : 
(2166,1084):(2230,1246) : 0
(2044,1084):(2166,1522) : 0
(1864,1400):(2044,1522) : 0
AN
use : z
dir : i
shape : 
(92,876):(274,1190) : 0
VSS
use : g
dir : b
shape : 
(2180,-160):(2800,160) : 0
(2000,-160):(2180,244) : 0
(1468,-160):(2000,160) : 0
(1288,-160):(1468,244) : 0
(612,-160):(1288,160) : 0
(432,-160):(612,244) : 0
(0,-160):(432,160) : 0
VDD
use : p
dir : b
shape : 
(2500,2240):(2800,2560) : 0
(2320,1942):(2500,2560) : 0
(670,2240):(2320,2560) : 0
(490,2130):(670,2560) : 0
(0,2240):(490,2560) : 0
NOR4BXL
--pins(7)
Y
use :  
dir : o
shape : 
(2072,878):(2080,988) : 0
(1944,574):(2072,1602) : 0
(1778,574):(1944,684) : 0
(1834,1440):(1944,1602) : 0
(856,522):(1778,684) : 0
D
use : 
dir : i
shape : 
(672,1112):(800,1510) : 0
(614,1400):(672,1510) : 0
(486,1400):(614,1522) : 0
C
use : 
dir : i
shape : 
(1056,1114):(1206,1276) : 0
(1016,878):(1056,1276) : 0
(928,878):(1016,1224) : 0
(852,878):(928,988) : 0
B
use :  
dir : i
shape : 
(1394,826):(1756,1026) : 0
AN
use : z
dir : i
shape : 
(76,790):(288,1064) : 0
VSS
use : g
dir : b
shape : 
(2088,-160):(2200,160) : 0
(1900,-160):(2088,244) : 0
(1356,-160):(1900,160) : 0
(1166,-160):(1356,244) : 0
(656,-160):(1166,160) : 0
(466,-160):(656,244) : 0
(0,-160):(466,160) : 0
VDD
use : p
dir : b
shape : 
(600,2240):(2200,2560) : 0
(412,2156):(600,2560) : 0
(0,2240):(412,2560) : 0
NOR4BX4
--pins(7)
Y
use :  
dir : o
shape : 
(6284,1134):(6324,1800) : 0
(6160,564):(6284,1846) : 0
(5816,564):(6160,674) : 0
(6120,1134):(6160,1846) : 0
(4786,1736):(6120,1846) : 0
(5632,512):(5816,674) : 0
(5032,564):(5632,674) : 0
(4848,512):(5032,674) : 0
(1832,564):(4848,674) : 0
(4728,1734):(4786,1896) : 0
(4604,1734):(4728,2016) : 0
(2060,1908):(4604,2016) : 0
(1878,1908):(2060,2070) : 0
(1648,512):(1832,674) : 0
(1056,564):(1648,674) : 0
(872,512):(1056,674) : 0
D
use : 
dir : i
shape : 
(5940,858):(6014,1020) : 0
(5816,858):(5940,1516) : 0
(3440,1408):(5816,1516) : 0
(3410,1408):(3440,1522) : 0
(3350,1236):(3410,1522) : 0
(3226,1236):(3350,1798) : 0
(818,1688):(3226,1798) : 0
(694,1052):(818,1798) : 0
C
use : 
dir : i
shape : 
(5578,952):(5638,1146) : 0
(5454,952):(5578,1296) : 0
(3890,1186):(5454,1296) : 0
(3766,1004):(3890,1296) : 0
(3706,1004):(3766,1166) : 0
(3630,1004):(3706,1146) : 0
(2958,1004):(3630,1114) : 0
(2898,1004):(2958,1166) : 0
(2770,1004):(2898,1578) : 0
(2604,1412):(2770,1578) : 0
(1210,1470):(2604,1578) : 0
(1056,1112):(1210,1578) : 0
(1026,1112):(1056,1274) : 0
B
use : 
dir : i
shape : 
(5094,914):(5276,1076) : 0
(4382,966):(5094,1076) : 0
(4234,866):(4382,1076) : 0
(4110,784):(4234,1076) : 0
(2554,784):(4110,892) : 0
(2430,784):(2554,1274) : 0
(2370,1112):(2430,1274) : 0
(1570,1146):(2370,1254) : 0
(1388,1126):(1570,1288) : 0
AN
use :  
dir : i
shape : 
(92,878):(274,1216) : 0
VSS
use : g
dir : b
shape : 
(6212,-160):(6400,160) : 0
(6028,-160):(6212,424) : 0
(5422,-160):(6028,160) : 0
(5240,-160):(5422,424) : 0
(4644,-160):(5240,160) : 0
(4460,-160):(4644,424) : 0
(2228,-160):(4460,160) : 0
(2044,-160):(2228,424) : 0
(1444,-160):(2044,160) : 0
(1260,-160):(1444,422) : 0
(668,-160):(1260,160) : 0
(484,-160):(668,422) : 0
(0,-160):(484,160) : 0
VDD
use : p
dir : b
shape : 
(6212,2240):(6400,2560) : 0
(6028,2156):(6212,2560) : 0
(3424,2240):(6028,2560) : 0
(3240,2156):(3424,2560) : 0
(698,2240):(3240,2560) : 0
(514,2156):(698,2560) : 0
(0,2240):(514,2560) : 0
NOR4BX2
--pins(7)
Y
use :  
dir : o
shape : 
(3350,384):(3474,1788) : 0
(3316,384):(3350,612) : 0
(2280,1678):(3350,1788) : 0
(1898,384):(3316,492) : 0
(2116,1666):(2280,1800) : 0
(1930,1652):(2116,1814) : 0
(1712,358):(1898,520) : 0
(884,384):(1712,492) : 0
D
use : 
dir : i
shape : 
(3160,1114):(3224,1276) : 0
(3038,1114):(3160,1522) : 0
(3036,1140):(3038,1522) : 0
(838,1412):(3036,1522) : 0
(780,1400):(838,1522) : 0
(594,1138):(780,1522) : 0
C
use :  
dir : i
shape : 
(2960,792):(3122,1000) : 0
(2800,686):(2960,1000) : 0
(1364,686):(2800,796) : 0
(1282,686):(1364,878) : 0
(1156,686):(1282,1066) : 0
B
use :  
dir : i
shape : 
(2278,904):(2552,1254) : 0
(1680,904):(2278,1014) : 0
(1494,904):(1680,1066) : 0
AN
use :  
dir : i
shape : 
(444,866):(644,1026) : 0
(320,790):(444,1026) : 0
VSS
use : g
dir : b
shape : 
(2312,-160):(3600,160) : 0
(2128,-160):(2312,244) : 0
(1484,-160):(2128,160) : 0
(1298,-160):(1484,244) : 0
(676,-160):(1298,160) : 0
(490,-160):(676,396) : 0
(0,-160):(490,160) : 0
VDD
use : p
dir : b
shape : 
(3448,2240):(3600,2560) : 0
(3262,2156):(3448,2560) : 0
(654,2240):(3262,2560) : 0
(470,2156):(654,2560) : 0
(0,2240):(470,2560) : 0
NOR4BX1
--pins(7)
Y
use :  
dir : o
shape : 
(2072,878):(2080,988) : 0
(1944,576):(2072,1598) : 0
(1778,576):(1944,686) : 0
(1834,1436):(1944,1598) : 0
(856,524):(1778,686) : 0
D
use : 
dir : i
shape : 
(672,1112):(800,1510) : 0
(614,1400):(672,1510) : 0
(486,1400):(614,1522) : 0
C
use :  
dir : i
shape : 
(1056,1114):(1206,1276) : 0
(1016,878):(1056,1276) : 0
(928,878):(1016,1224) : 0
(852,878):(928,988) : 0
B
use :  
dir : i
shape : 
(1394,826):(1756,1026) : 0
AN
use :  
dir : i
shape : 
(286,790):(288,1062) : 0
(98,790):(286,1064) : 0
(76,790):(98,1062) : 0
VSS
use : g
dir : b
shape : 
(2088,-160):(2200,160) : 0
(1900,-160):(2088,244) : 0
(1356,-160):(1900,160) : 0
(1166,-160):(1356,244) : 0
(656,-160):(1166,160) : 0
(466,-160):(656,244) : 0
(0,-160):(466,160) : 0
VDD
use : p
dir : b
shape : 
(656,2240):(2200,2560) : 0
(466,2156):(656,2560) : 0
(0,2240):(466,2560) : 0
NOR4X2
--pins(7)
Y
use :  
dir : o
shape : 
(2960,574):(3084,2016) : 0
(1626,574):(2960,684) : 0
(2920,1788):(2960,2016) : 0
(1706,1908):(2920,2016) : 0
(1522,1908):(1706,2070) : 0
(1444,522):(1626,684) : 0
(676,574):(1444,684) : 0
(492,522):(676,684) : 0
D
use : 
dir : i
shape : 
(2774,1112):(2834,1274) : 0
(2650,1112):(2774,1798) : 0
(476,1688):(2650,1798) : 0
(352,1112):(476,1798) : 0
(110,1112):(352,1274) : 0
C
use :  
dir : i
shape : 
(2348,792):(2472,1578) : 0
(2290,792):(2348,954) : 0
(950,1470):(2348,1578) : 0
(854,1412):(950,1578) : 0
(730,1112):(854,1578) : 0
(670,1112):(730,1274) : 0
B
use :  
dir : i
shape : 
(2138,1112):(2198,1274) : 0
(2014,888):(2138,1274) : 0
(1306,888):(2014,998) : 0
(1214,878):(1306,998) : 0
(1034,878):(1214,1076) : 0
(1032,914):(1034,1076) : 0
A
use :  
dir : i
shape : 
(1420,1110):(1756,1272) : 0
VSS
use : g
dir : b
shape : 
(2036,-160):(3200,160) : 0
(1854,-160):(2036,244) : 0
(1186,-160):(1854,160) : 0
(1002,-160):(1186,244) : 0
(280,-160):(1002,160) : 0
(96,-160):(280,450) : 0
(0,-160):(96,160) : 0
VDD
use : p
dir : b
shape : 
(3068,2240):(3200,2560) : 0
(2884,2156):(3068,2560) : 0
(280,2240):(2884,2560) : 0
(96,2156):(280,2560) : 0
(0,2240):(96,2560) : 0
NOR4X1
--pins(7)
Y
use :  
dir : o
shape : 
(1952,538):(2080,1522) : 0
(522,538):(1952,700) : 0
(1758,1412):(1952,1522) : 0
(1570,1396):(1758,1780) : 0
D
use : 
dir : i
shape : 
(312,1084):(314,1246) : 0
(124,1084):(312,1400) : 0
(114,1146):(124,1254) : 0
C
use :  
dir : i
shape : 
(486,842):(880,1038) : 0
B
use :  
dir : i
shape : 
(1186,866):(1252,1028) : 0
(1058,866):(1186,1522) : 0
(852,1400):(1058,1522) : 0
A
use :  
dir : i
shape : 
(1622,840):(1812,1120) : 0
(1586,878):(1622,988) : 0
VSS
use : g
dir : b
shape : 
(2100,-160):(2200,160) : 0
(1912,-160):(2100,244) : 0
(1222,-160):(1912,160) : 0
(1034,-160):(1222,244) : 0
(288,-160):(1034,160) : 0
(100,-160):(288,244) : 0
(0,-160):(100,160) : 0
VDD
use : p
dir : b
shape : 
(288,2240):(2200,2560) : 0
(100,2156):(288,2560) : 0
(0,2240):(100,2560) : 0
NOR3BX4
--pins(6)
Y
use :  
dir : o
shape : 
(3840,866):(3922,1704) : 0
(3714,536):(3840,1704) : 0
(2862,536):(3714,646) : 0
(3614,1542):(3714,1704) : 0
(2104,1542):(3614,1652) : 0
(2736,330):(2862,646) : 0
(2674,330):(2736,492) : 0
(2022,384):(2674,492) : 0
(2064,1542):(2104,1678) : 0
(1936,1542):(2064,1734) : 0
(1834,330):(2022,492) : 0
(1752,1624):(1936,1734) : 0
(1184,384):(1834,492) : 0
(1564,1624):(1752,1786) : 0
(998,330):(1184,492) : 0
C
use : 
dir : i
shape : 
(2590,828):(2910,990) : 0
(2462,602):(2590,990) : 0
(972,602):(2462,712) : 0
(846,602):(972,1254) : 0
(732,1072):(846,1234) : 0
B
use :  
dir : i
shape : 
(3122,1046):(3248,1212) : 0
(2256,1102):(3122,1212) : 0
(2196,1040):(2256,1212) : 0
(2068,822):(2196,1212) : 0
(2064,822):(2068,1000) : 0
(1336,822):(2064,930) : 0
(1316,822):(1336,1026) : 0
(1130,822):(1316,1028) : 0
AN
use :  
dir : i
shape : 
(568,612):(608,722) : 0
(440,612):(568,1038) : 0
(360,876):(440,1038) : 0
VSS
use : g
dir : b
shape : 
(3258,-160):(4000,160) : 0
(3072,-160):(3258,396) : 0
(2444,-160):(3072,160) : 0
(2256,-160):(2444,244) : 0
(1604,-160):(2256,160) : 0
(1416,-160):(1604,244) : 0
(788,-160):(1416,160) : 0
(600,-160):(788,396) : 0
(0,-160):(600,160) : 0
VDD
use : p
dir : b
shape : 
(2776,2240):(4000,2560) : 0
(2590,1822):(2776,2560) : 0
(716,2240):(2590,2560) : 0
(528,1732):(716,2560) : 0
(0,2240):(528,2560) : 0
NOR3BX2
--pins(6)
Y
use :  
dir : o
shape : 
(2540,384):(2662,1722) : 0
(2524,384):(2540,612) : 0
(2524,1522):(2540,1722) : 0
(1946,384):(2524,492) : 0
(1986,1612):(2524,1722) : 0
(1864,1612):(1986,1788) : 0
(1766,330):(1946,492) : 0
(1686,1612):(1864,1722) : 0
(1140,384):(1766,492) : 0
(1506,1612):(1686,1790) : 0
(960,330):(1140,492) : 0
C
use : 
dir : i
shape : 
(2360,788):(2418,950) : 0
(2238,648):(2360,950) : 0
(934,648):(2238,758) : 0
(934,1146):(936,1254) : 0
(812,648):(934,1254) : 0
(774,988):(812,1254) : 0
(730,1072):(774,1254) : 0
(670,1072):(730,1234) : 0
B
use :  
dir : i
shape : 
(2114,1110):(2172,1272) : 0
(1992,922):(2114,1272) : 0
(1286,922):(1992,1030) : 0
(1238,878):(1286,1030) : 0
(1116,878):(1238,1084) : 0
AN
use :  
dir : i
shape : 
(546,612):(586,722) : 0
(424,612):(546,914) : 0
(348,752):(424,914) : 0
VSS
use : g
dir : b
shape : 
(1544,-160):(2800,160) : 0
(1362,-160):(1544,244) : 0
(758,-160):(1362,160) : 0
(578,-160):(758,396) : 0
(0,-160):(578,160) : 0
VDD
use : p
dir : b
shape : 
(2672,2240):(2800,2560) : 0
(2492,1864):(2672,2560) : 0
(690,2240):(2492,2560) : 0
(510,1794):(690,2560) : 0
(0,2240):(510,2560) : 0
NOR3BX1
--pins(6)
Y
use :  
dir : o
shape : 
(2006,538):(2134,1788) : 0
(972,538):(2006,700) : 0
(1756,1678):(2006,1788) : 0
(1566,1678):(1756,1848) : 0
C
use : 
dir : i
shape : 
(978,1146):(980,1254) : 0
(614,1072):(978,1254) : 0
B
use :  
dir : i
shape : 
(1106,828):(1512,1022) : 0
AN
use :  
dir : i
shape : 
(572,612):(614,722) : 0
(444,612):(572,914) : 0
(364,752):(444,914) : 0
VSS
use : g
dir : b
shape : 
(1584,-160):(2200,160) : 0
(1394,-160):(1584,244) : 0
(830,-160):(1394,160) : 0
(642,-160):(830,244) : 0
(0,-160):(642,160) : 0
VDD
use : p
dir : b
shape : 
(722,2240):(2200,2560) : 0
(534,1794):(722,2560) : 0
(0,2240):(534,2560) : 0
NOR3X4
--pins(6)
Y
use :  
dir : o
shape : 
(3442,1134):(3524,1800) : 0
(3316,536):(3442,1800) : 0
(2248,536):(3316,646) : 0
(3122,1620):(3316,1784) : 0
(1330,1674):(3122,1784) : 0
(2062,484):(2248,646) : 0
(1462,536):(2062,646) : 0
(1276,484):(1462,646) : 0
(1146,1674):(1330,1836) : 0
(676,536):(1276,646) : 0
(490,484):(676,646) : 0
C
use : 
dir : i
shape : 
(2184,1196):(2378,1548) : 0
(2042,1400):(2184,1548) : 0
(306,1438):(2042,1548) : 0
(180,1052):(306,1548) : 0
(112,1052):(180,1254) : 0
B
use :  
dir : i
shape : 
(1942,976):(2780,1086) : 0
(1816,976):(1942,1220) : 0
(808,1110):(1816,1220) : 0
(748,1014):(808,1220) : 0
(622,878):(748,1220) : 0
(478,878):(622,988) : 0
A
use :  
dir : i
shape : 
(3106,1162):(3164,1324) : 0
(2980,758):(3106,1324) : 0
(1462,758):(2980,866) : 0
(2978,1162):(2980,1324) : 0
(1276,758):(1462,992) : 0
(1198,858):(1276,988) : 0
VSS
use : g
dir : b
shape : 
(2640,-160):(3600,160) : 0
(2454,-160):(2640,396) : 0
(1854,-160):(2454,160) : 0
(1670,-160):(1854,396) : 0
(1070,-160):(1670,160) : 0
(884,-160):(1070,396) : 0
(284,-160):(884,160) : 0
(98,-160):(284,422) : 0
(0,-160):(98,160) : 0
VDD
use : p
dir : b
shape : 
(2362,2240):(3600,2560) : 0
(2176,1978):(2362,2560) : 0
(284,2240):(2176,2560) : 0
(98,1858):(284,2560) : 0
(0,2240):(98,2560) : 0
NOR3X2
--pins(6)
Y
use :  
dir : o
shape : 
(2350,510):(2480,1710) : 0
(1508,510):(2350,620) : 0
(2308,1534):(2350,1710) : 0
(1374,1600):(2308,1710) : 0
(1316,302):(1508,688) : 0
(1182,1600):(1374,1780) : 0
(698,578):(1316,688) : 0
(506,302):(698,688) : 0
C
use : 
dir : i
shape : 
(2014,1074):(2176,1488) : 0
(428,1378):(2014,1488) : 0
(298,1146):(428,1488) : 0
(236,1146):(298,1414) : 0
(116,1146):(236,1254) : 0
B
use :  
dir : i
shape : 
(1826,754):(1886,916) : 0
(1696,754):(1826,1270) : 0
(1694,754):(1696,916) : 0
(832,1160):(1696,1270) : 0
(830,916):(832,1270) : 0
(704,890):(830,1270) : 0
(642,890):(704,1078) : 0
(622,890):(642,1000) : 0
(492,878):(622,1000) : 0
A
use :  
dir : i
shape : 
(996,878):(1364,1050) : 0
VSS
use : g
dir : b
shape : 
(1104,-160):(2600,160) : 0
(912,-160):(1104,422) : 0
(292,-160):(912,160) : 0
(102,-160):(292,422) : 0
(0,-160):(102,160) : 0
VDD
use : p
dir : b
shape : 
(2408,2240):(2600,2560) : 0
(2218,1850):(2408,2560) : 0
(292,2240):(2218,2560) : 0
(102,1752):(292,2560) : 0
(0,2240):(102,2560) : 0
NOR3X1
--pins(6)
Y
use :  
dir : o
shape : 
(1332,538):(1336,1788) : 0
(1214,538):(1332,1848) : 0
(392,538):(1214,700) : 0
(1114,1678):(1214,1848) : 0
C
use : 
dir : i
shape : 
(274,1072):(276,1234) : 0
(96,1072):(274,1388) : 0
B
use :  
dir : i
shape : 
(464,842):(722,1122) : 0
A
use :  
dir : i
shape : 
(1034,1072):(1092,1234) : 0
(912,1072):(1034,1522) : 0
(814,1412):(912,1522) : 0
VSS
use : g
dir : b
shape : 
(870,-160):(1400,160) : 0
(690,-160):(870,244) : 0
(276,-160):(690,160) : 0
(96,-160):(276,244) : 0
(0,-160):(96,160) : 0
VDD
use : p
dir : b
shape : 
(276,2240):(1400,2560) : 0
(96,1800):(276,2560) : 0
(0,2240):(96,2560) : 0
NOR2BXL
--pins(5)
Y
use :  
dir : o
shape : 
(1210,590):(1332,1596) : 0
(1002,590):(1210,700) : 0
(1124,1412):(1210,1596) : 0
(822,538):(1002,700) : 0
B
use : 
dir : i
shape : 
(822,1134):(1050,1266) : 0
(642,1134):(822,1324) : 0
AN
use :  
dir : i
shape : 
(74,866):(276,1162) : 0
VSS
use : g
dir : b
shape : 
(1304,-160):(1400,160) : 0
(1124,-160):(1304,244) : 0
(626,-160):(1124,160) : 0
(446,-160):(626,244) : 0
(0,-160):(446,160) : 0
VDD
use : p
dir : b
shape : 
(604,2240):(1400,2560) : 0
(424,2156):(604,2560) : 0
(0,2240):(424,2560) : 0
NOR2BX4
--pins(5)
Y
use :  
dir : o
shape : 
(2524,528):(2726,1572) : 0
(1946,528):(2524,672) : 0
(2504,1386):(2524,1572) : 0
(1146,1410):(2504,1572) : 0
(1766,510):(1946,672) : 0
(1140,562):(1766,672) : 0
(960,510):(1140,672) : 0
B
use : 
dir : i
shape : 
(1872,1126):(2052,1300) : 0
(936,1190):(1872,1300) : 0
(822,1130):(936,1300) : 0
(642,1042):(822,1300) : 0
AN
use :  
dir : i
shape : 
(68,872):(276,1142) : 0
VSS
use : g
dir : b
shape : 
(2354,-160):(2800,160) : 0
(2174,-160):(2354,244) : 0
(1544,-160):(2174,160) : 0
(1362,-160):(1544,244) : 0
(732,-160):(1362,160) : 0
(552,-160):(732,244) : 0
(0,-160):(552,160) : 0
VDD
use : p
dir : b
shape : 
(2026,2240):(2800,2560) : 0
(1846,2156):(2026,2560) : 0
(626,2234):(1846,2560) : 0
(446,2156):(626,2560) : 0
(0,2240):(446,2560) : 0
NOR2BX2
--pins(5)
Y
use :  
dir : o
shape : 
(1994,616):(2122,1534) : 0
(1700,616):(1994,726) : 0
(1952,1412):(1994,1534) : 0
(1378,1424):(1952,1534) : 0
(1512,564):(1700,726) : 0
(1188,1424):(1378,1586) : 0
B
use : 
dir : i
shape : 
(1694,836):(1856,1130) : 0
(1022,836):(1694,946) : 0
(872,600):(1022,946) : 0
(812,600):(872,1028) : 0
(714,836):(812,1028) : 0
(684,866):(714,1028) : 0
AN
use :  
dir : i
shape : 
(100,914):(288,1266) : 0
VSS
use : g
dir : b
shape : 
(2100,-160):(2200,160) : 0
(1912,-160):(2100,456) : 0
(1272,-160):(1912,160) : 0
(1084,-160):(1272,244) : 0
(0,-160):(1084,160) : 0
VDD
use : p
dir : b
shape : 
(2100,2240):(2200,2560) : 0
(1912,2156):(2100,2560) : 0
(644,2240):(1912,2560) : 0
(456,2156):(644,2560) : 0
(0,2240):(456,2560) : 0
NOR2BX1
--pins(5)
Y
use :  
dir : o
shape : 
(1210,590):(1332,1716) : 0
(1002,590):(1210,700) : 0
(1124,1412):(1210,1716) : 0
(822,538):(1002,700) : 0
B
use : 
dir : i
shape : 
(822,1134):(1050,1266) : 0
(642,1134):(822,1340) : 0
AN
use :  
dir : i
shape : 
(74,972):(276,1266) : 0
VSS
use : g
dir : b
shape : 
(1304,-160):(1400,160) : 0
(1124,-160):(1304,244) : 0
(706,-160):(1124,160) : 0
(526,-160):(706,244) : 0
(0,-160):(526,160) : 0
VDD
use : p
dir : b
shape : 
(604,2240):(1400,2560) : 0
(424,1832):(604,2560) : 0
(0,2240):(424,2560) : 0
NOR2XL
--pins(5)
Y
use :  
dir : o
shape : 
(982,590):(1122,1548) : 0
(704,590):(982,700) : 0
(884,1252):(982,1548) : 0
(496,538):(704,700) : 0
B
use : 
dir : i
shape : 
(328,1134):(510,1266) : 0
(122,1096):(328,1266) : 0
(84,1134):(122,1266) : 0
A
use :  
dir : i
shape : 
(484,812):(842,1004) : 0
VSS
use : g
dir : b
shape : 
(1090,-160):(1200,160) : 0
(884,-160):(1090,244) : 0
(316,-160):(884,160) : 0
(110,-160):(316,244) : 0
(0,-160):(110,160) : 0
VDD
use : p
dir : b
shape : 
(316,2240):(1200,2560) : 0
(110,2156):(316,2560) : 0
(0,2240):(110,2560) : 0
NOR2X4
--pins(5)
Y
use :  
dir : o
shape : 
(2498,866):(2522,1534) : 0
(2488,530):(2498,1534) : 0
(2330,530):(2488,1680) : 0
(1530,530):(2330,674) : 0
(2308,866):(2330,1680) : 0
(2296,1386):(2308,1680) : 0
(856,1520):(2296,1680) : 0
(1340,512):(1530,674) : 0
(720,564):(1340,674) : 0
(530,512):(720,674) : 0
B
use : 
dir : i
shape : 
(1654,1122):(1716,1284) : 0
(1526,1122):(1654,1410) : 0
(622,1300):(1526,1410) : 0
(492,1300):(622,1522) : 0
(468,1300):(492,1414) : 0
(338,984):(468,1414) : 0
(276,984):(338,1146) : 0
A
use :  
dir : i
shape : 
(2110,928):(2172,1090) : 0
(1980,788):(2110,1090) : 0
(1046,788):(1980,898) : 0
(918,788):(1046,1050) : 0
(864,878):(918,1050) : 0
(856,940):(864,1050) : 0
VSS
use : g
dir : b
shape : 
(1958,-160):(2600,160) : 0
(1768,-160):(1958,244) : 0
(1126,-160):(1768,160) : 0
(934,-160):(1126,422) : 0
(292,-160):(934,160) : 0
(102,-160):(292,596) : 0
(0,-160):(102,160) : 0
VDD
use : p
dir : b
shape : 
(1790,2240):(2600,2560) : 0
(1598,2156):(1790,2560) : 0
(304,2240):(1598,2560) : 0
(112,2156):(304,2560) : 0
(0,2240):(112,2560) : 0
NOR2X2
--pins(5)
Y
use :  
dir : o
shape : 
(1724,616):(1734,1522) : 0
(1610,616):(1724,1534) : 0
(1310,616):(1610,726) : 0
(1558,1412):(1610,1534) : 0
(992,1424):(1558,1534) : 0
(1124,340):(1310,726) : 0
(808,1424):(992,1586) : 0
B
use : 
dir : i
shape : 
(1304,836):(1484,1128) : 0
(458,836):(1304,946) : 0
(240,836):(458,1036) : 0
(118,836):(240,988) : 0
A
use :  
dir : i
shape : 
(654,1076):(1004,1266) : 0
VSS
use : g
dir : b
shape : 
(1702,-160):(1800,160) : 0
(1516,-160):(1702,456) : 0
(916,-160):(1516,160) : 0
(730,-160):(916,680) : 0
(0,-160):(730,160) : 0
VDD
use : p
dir : b
shape : 
(1702,2240):(1800,2560) : 0
(1516,2156):(1702,2560) : 0
(284,2240):(1516,2560) : 0
(98,2156):(284,2560) : 0
(0,2240):(98,2560) : 0
NOR2X1
--pins(5)
Y
use :  
dir : o
shape : 
(982,590):(1122,1548) : 0
(704,590):(982,700) : 0
(884,1252):(982,1548) : 0
(496,538):(704,700) : 0
B
use : 
dir : i
shape : 
(328,1134):(510,1286) : 0
(122,1096):(328,1286) : 0
(84,1134):(122,1286) : 0
A
use :  
dir : i
shape : 
(484,814):(842,1004) : 0
VSS
use : g
dir : b
shape : 
(1090,-160):(1200,160) : 0
(884,-160):(1090,244) : 0
(316,-160):(884,160) : 0
(110,-160):(316,244) : 0
(0,-160):(110,160) : 0
VDD
use : p
dir : b
shape : 
(316,2240):(1200,2560) : 0
(110,2156):(316,2560) : 0
(0,2240):(110,2560) : 0
NAND4BBX1
--pins(7)
Y
use :  
dir : o
shape : 
(2686,1146):(2734,1866) : 0
(2612,402):(2686,1866) : 0
(2564,402):(2612,1254) : 0
(1756,1758):(2612,1866) : 0
(2524,402):(2564,612) : 0
(1928,402):(2524,512) : 0
(1748,402):(1928,564) : 0
(1634,1484):(1756,1866) : 0
(1576,1484):(1634,1678) : 0
(1474,1510):(1576,1678) : 0
(1164,1510):(1474,1620) : 0
(1034,1484):(1164,1620) : 0
(854,1484):(1034,1646) : 0
D
use : 
dir : i
shape : 
(824,878):(936,988) : 0
(702,878):(824,1200) : 0
(654,1038):(702,1200) : 0
C
use :  
dir : i
shape : 
(1220,878):(1286,988) : 0
(1098,878):(1220,1272) : 0
(1004,1110):(1098,1272) : 0
BN
use :  
dir : i
shape : 
(82,866):(284,1148) : 0
AN
use :  
dir : i
shape : 
(2376,996):(2402,1158) : 0
(2140,996):(2376,1266) : 0
VSS
use : g
dir : b
shape : 
(2704,-160):(2800,160) : 0
(2524,-160):(2704,244) : 0
(632,-160):(2524,160) : 0
(196,-160):(632,244) : 0
(0,-160):(196,160) : 0
VDD
use : p
dir : b
shape : 
(2154,2240):(2800,2560) : 0
(1914,2156):(2154,2560) : 0
(1394,2240):(1914,2560) : 0
(1214,2156):(1394,2560) : 0
(674,2240):(1214,2560) : 0
(644,2156):(674,2560) : 0
(522,2130):(644,2560) : 0
(494,2156):(522,2560) : 0
(0,2240):(494,2560) : 0
NAND4BXL
--pins(7)
Y
use :  
dir : o
shape : 
(1336,1678):(1714,1788) : 0
(1344,504):(1534,666) : 0
(1278,558):(1344,666) : 0
(1278,1678):(1336,1878) : 0
(1150,558):(1278,1878) : 0
(980,1716):(1150,1878) : 0
(600,1770):(980,1878) : 0
(412,1716):(600,1878) : 0
D
use : 
dir : i
shape : 
(156,878):(334,1200) : 0
(120,878):(156,1198) : 0
C
use :  
dir : i
shape : 
(444,1322):(766,1534) : 0
B
use :  
dir : i
shape : 
(736,866):(1022,1064) : 0
AN
use :  
dir : i
shape : 
(1748,1092):(2122,1304) : 0
VSS
use : g
dir : b
shape : 
(1914,-160):(2200,160) : 0
(1726,-160):(1914,244) : 0
(288,-160):(1726,160) : 0
(100,-160):(288,244) : 0
(0,-160):(100,160) : 0
VDD
use : p
dir : b
shape : 
(1764,2240):(2200,2560) : 0
(1574,2156):(1764,2560) : 0
(1022,2240):(1574,2560) : 0
(834,2156):(1022,2560) : 0
(288,2240):(834,2560) : 0
(100,2156):(288,2560) : 0
(0,2240):(100,2560) : 0
NAND4BX4
--pins(7)
Y
use :  
dir : o
shape : 
(5966,1134):(5970,1800) : 0
(5948,576):(5966,1800) : 0
(5842,576):(5948,1884) : 0
(4632,576):(5842,686) : 0
(5764,1134):(5842,1884) : 0
(4588,1740):(5764,1884) : 0
(4450,300):(4632,686) : 0
(934,1740):(4588,1874) : 0
(2004,414):(4450,548) : 0
(1820,300):(2004,686) : 0
D
use : 
dir : i
shape : 
(5630,852):(5718,1014) : 0
(5538,852):(5630,1630) : 0
(5506,878):(5538,1630) : 0
(3318,1522):(5506,1630) : 0
(3136,1470):(3318,1630) : 0
(950,1522):(3136,1630) : 0
(906,1412):(950,1630) : 0
(826,1038):(906,1630) : 0
(782,1038):(826,1522) : 0
(722,1038):(782,1200) : 0
C
use :  
dir : i
shape : 
(5336,1038):(5366,1200) : 0
(5182,1038):(5336,1266) : 0
(5178,1146):(5182,1266) : 0
(5094,1146):(5178,1412) : 0
(5054,1158):(5094,1412) : 0
(3832,1302):(5054,1412) : 0
(3650,1250):(3832,1412) : 0
(2802,1250):(3650,1360) : 0
(2618,1250):(2802,1412) : 0
(1306,1302):(2618,1412) : 0
(1182,1038):(1306,1412) : 0
(1088,1038):(1182,1200) : 0
B
use :  
dir : i
shape : 
(4902,1030):(4930,1192) : 0
(4698,866):(4902,1192) : 0
(4208,1084):(4698,1192) : 0
(4006,1020):(4208,1192) : 0
(2444,1020):(4006,1128) : 0
(2242,1020):(2444,1192) : 0
(1648,1084):(2242,1192) : 0
(1446,1030):(1648,1192) : 0
AN
use :  
dir : i
shape : 
(84,866):(288,1148) : 0
VSS
use : g
dir : b
shape : 
(5948,-160):(6400,160) : 0
(5764,-160):(5948,244) : 0
(3318,-160):(5764,160) : 0
(3136,-160):(3318,244) : 0
(690,-160):(3136,160) : 0
(506,-160):(690,244) : 0
(0,-160):(506,160) : 0
VDD
use : p
dir : b
shape : 
(5902,2240):(6400,2560) : 0
(5718,2156):(5902,2560) : 0
(5136,2240):(5718,2560) : 0
(4954,2156):(5136,2560) : 0
(4398,2240):(4954,2560) : 0
(4156,2156):(4398,2560) : 0
(2298,2240):(4156,2560) : 0
(2056,2156):(2298,2560) : 0
(1500,2240):(2056,2560) : 0
(1318,2156):(1500,2560) : 0
(736,2240):(1318,2560) : 0
(552,2156):(736,2560) : 0
(0,2240):(552,2560) : 0
NAND4BX2
--pins(7)
Y
use :  
dir : o
shape : 
(3480,390):(3482,1266) : 0
(3330,390):(3480,1946) : 0
(3316,390):(3330,612) : 0
(3316,1128):(3330,1946) : 0
(1974,390):(3316,524) : 0
(2090,1802):(3316,1946) : 0
(1926,1740):(2090,1946) : 0
(1790,300):(1974,686) : 0
(878,1740):(1926,1884) : 0
D
use : 
dir : i
shape : 
(2714,1522):(2900,1684) : 0
(962,1522):(2714,1630) : 0
(848,1412):(962,1630) : 0
(838,1038):(848,1630) : 0
(722,1038):(838,1522) : 0
(680,1038):(722,1200) : 0
C
use :  
dir : i
shape : 
(2754,1146):(2762,1254) : 0
(2694,1038):(2754,1254) : 0
(2570,1038):(2694,1412) : 0
(1254,1302):(2570,1412) : 0
(1130,1038):(1254,1412) : 0
(1042,1038):(1130,1200) : 0
B
use :  
dir : i
shape : 
(2376,878):(2402,988) : 0
(2236,866):(2376,1192) : 0
(2170,1028):(2236,1192) : 0
(1600,1084):(2170,1192) : 0
(1396,1030):(1600,1192) : 0
AN
use :  
dir : i
shape : 
(84,866):(292,1148) : 0
VSS
use : g
dir : b
shape : 
(3306,-160):(3600,160) : 0
(3120,-160):(3306,244) : 0
(644,-160):(3120,160) : 0
(458,-160):(644,244) : 0
(0,-160):(458,160) : 0
VDD
use : p
dir : b
shape : 
(2258,2240):(3600,2560) : 0
(2012,2156):(2258,2560) : 0
(1450,2240):(2012,2560) : 0
(1266,2156):(1450,2560) : 0
(676,2240):(1266,2560) : 0
(646,2156):(676,2560) : 0
(520,2130):(646,2560) : 0
(490,2156):(520,2560) : 0
(0,2240):(490,2560) : 0
NAND4BX1
--pins(7)
Y
use :  
dir : o
shape : 
(2480,1146):(2530,1866) : 0
(2400,402):(2480,1866) : 0
(2350,402):(2400,1254) : 0
(1492,1758):(2400,1866) : 0
(2308,402):(2350,612) : 0
(1674,402):(2308,512) : 0
(1482,402):(1674,564) : 0
(1362,1474):(1492,1866) : 0
(1300,1474):(1362,1678) : 0
(1194,1526):(1300,1678) : 0
(726,1526):(1194,1636) : 0
(534,1474):(726,1636) : 0
D
use : 
dir : i
shape : 
(504,878):(622,988) : 0
(374,878):(504,1200) : 0
(324,984):(374,1200) : 0
C
use :  
dir : i
shape : 
(932,878):(994,988) : 0
(886,878):(932,1246) : 0
(802,878):(886,1272) : 0
(696,1110):(802,1272) : 0
B
use :  
dir : i
shape : 
(1134,1110):(1486,1330) : 0
AN
use :  
dir : i
shape : 
(2150,996):(2178,1158) : 0
(1900,996):(2150,1266) : 0
VSS
use : g
dir : b
shape : 
(2498,-160):(2600,160) : 0
(2308,-160):(2498,244) : 0
(302,-160):(2308,160) : 0
(110,-160):(302,244) : 0
(0,-160):(110,160) : 0
VDD
use : p
dir : b
shape : 
(1914,2240):(2600,2560) : 0
(1660,2156):(1914,2560) : 0
(1108,2240):(1660,2560) : 0
(918,2156):(1108,2560) : 0
(348,2240):(918,2560) : 0
(158,2156):(348,2560) : 0
(0,2240):(158,2560) : 0
NAND4XL
--pins(7)
Y
use :  
dir : o
shape : 
(1320,592):(1622,754) : 0
(1184,1474):(1370,1636) : 0
(962,646):(1320,754) : 0
(962,1474):(1184,1584) : 0
(838,646):(962,1584) : 0
(616,1474):(838,1584) : 0
(430,1474):(616,1636) : 0
D
use : 
dir : i
shape : 
(284,1116):(352,1278) : 0
(158,878):(284,1278) : 0
(118,878):(158,988) : 0
C
use :  
dir : i
shape : 
(660,1116):(692,1278) : 0
(534,878):(660,1278) : 0
(478,878):(534,988) : 0
B
use :  
dir : i
shape : 
(1246,878):(1322,988) : 0
(1120,878):(1246,1278) : 0
(1088,1116):(1120,1278) : 0
A
use :  
dir : i
shape : 
(1674,878):(1682,988) : 0
(1516,878):(1674,1278) : 0
(1490,1116):(1516,1278) : 0
VSS
use : g
dir : b
shape : 
(292,-160):(1800,160) : 0
(106,-160):(292,244) : 0
(0,-160):(106,160) : 0
VDD
use : p
dir : b
shape : 
(1702,2240):(1800,2560) : 0
(1516,2156):(1702,2560) : 0
(1138,2240):(1516,2560) : 0
(944,2156):(1138,2560) : 0
(284,2240):(944,2560) : 0
(98,2156):(284,2560) : 0
(0,2240):(98,2560) : 0
NAND4X4
--pins(7)
Y
use :  
dir : o
shape : 
(5572,384):(5606,1278) : 0
(5550,384):(5572,1800) : 0
(5446,384):(5550,1884) : 0
(5368,384):(5446,614) : 0
(5368,1134):(5446,1884) : 0
(4352,384):(5368,526) : 0
(4200,1740):(5368,1884) : 0
(4246,300):(4352,526) : 0
(4064,300):(4246,686) : 0
(574,1740):(4200,1874) : 0
(1636,414):(4064,548) : 0
(1454,300):(1636,686) : 0
D
use : 
dir : i
shape : 
(5236,852):(5324,1014) : 0
(5144,852):(5236,1630) : 0
(5112,878):(5144,1630) : 0
(2942,1522):(5112,1630) : 0
(2760,1470):(2942,1630) : 0
(590,1522):(2760,1630) : 0
(546,1412):(590,1630) : 0
(468,1038):(546,1630) : 0
(422,1038):(468,1522) : 0
(364,1038):(422,1200) : 0
C
use :  
dir : i
shape : 
(4944,1038):(4974,1200) : 0
(4792,1038):(4944,1266) : 0
(4786,1146):(4792,1266) : 0
(4704,1146):(4786,1412) : 0
(4664,1158):(4704,1412) : 0
(3452,1302):(4664,1412) : 0
(3270,1250):(3452,1412) : 0
(2428,1250):(3270,1360) : 0
(2246,1250):(2428,1412) : 0
(944,1302):(2246,1412) : 0
(820,1038):(944,1412) : 0
(728,1038):(820,1200) : 0
B
use :  
dir : i
shape : 
(4514,1030):(4540,1192) : 0
(4310,866):(4514,1192) : 0
(3824,1084):(4310,1192) : 0
(3622,1020):(3824,1192) : 0
(2072,1020):(3622,1128) : 0
(1872,1020):(2072,1192) : 0
(1284,1084):(1872,1192) : 0
(1082,1030):(1284,1192) : 0
A
use :  
dir : i
shape : 
(3976,800):(4176,974) : 0
(1652,800):(3976,910) : 0
(1452,800):(1652,974) : 0
(984,800):(1452,910) : 0
(860,612):(984,910) : 0
(820,612):(860,722) : 0
VSS
use : g
dir : b
shape : 
(5550,-160):(6000,160) : 0
(5368,-160):(5550,244) : 0
(2942,-160):(5368,160) : 0
(2760,-160):(2942,244) : 0
(332,-160):(2760,160) : 0
(150,-160):(332,244) : 0
(0,-160):(150,160) : 0
VDD
use : p
dir : b
shape : 
(5506,2240):(6000,2560) : 0
(5324,2156):(5506,2560) : 0
(4746,2240):(5324,2560) : 0
(4564,2156):(4746,2560) : 0
(4014,2240):(4564,2560) : 0
(3772,2156):(4014,2560) : 0
(1928,2240):(3772,2560) : 0
(1688,2156):(1928,2560) : 0
(1136,2240):(1688,2560) : 0
(954,2156):(1136,2560) : 0
(378,2240):(954,2560) : 0
(196,2156):(378,2560) : 0
(0,2240):(196,2560) : 0
NAND4X2
--pins(7)
Y
use :  
dir : o
shape : 
(3082,390):(3084,1266) : 0
(2934,390):(3082,1946) : 0
(2920,390):(2934,612) : 0
(2920,1128):(2934,1946) : 0
(1594,390):(2920,524) : 0
(1708,1802):(2920,1946) : 0
(1546,1740):(1708,1946) : 0
(1412,300):(1594,686) : 0
(512,1740):(1546,1884) : 0
D
use : 
dir : i
shape : 
(2324,1522):(2508,1684) : 0
(596,1522):(2324,1630) : 0
(482,1412):(596,1630) : 0
(472,1038):(482,1630) : 0
(358,1038):(472,1522) : 0
(298,1038):(358,1200) : 0
C
use :  
dir : i
shape : 
(2374,1038):(2386,1200) : 0
(2328,1038):(2374,1254) : 0
(2204,1038):(2328,1412) : 0
(884,1302):(2204,1412) : 0
(760,1038):(884,1412) : 0
(666,1038):(760,1200) : 0
B
use :  
dir : i
shape : 
(1832,878):(2034,1192) : 0
(1226,1084):(1832,1192) : 0
(1024,1030):(1226,1192) : 0
A
use :  
dir : i
shape : 
(1396,802):(1598,974) : 0
(992,802):(1396,912) : 0
(868,612):(992,912) : 0
(826,612):(868,722) : 0
VSS
use : g
dir : b
shape : 
(2910,-160):(3200,160) : 0
(2726,-160):(2910,244) : 0
(280,-160):(2726,160) : 0
(96,-160):(280,244) : 0
(0,-160):(96,160) : 0
VDD
use : p
dir : b
shape : 
(1874,2240):(3200,2560) : 0
(1632,2156):(1874,2560) : 0
(1078,2240):(1632,2560) : 0
(894,2156):(1078,2560) : 0
(312,2240):(894,2560) : 0
(130,2156):(312,2560) : 0
(0,2240):(130,2560) : 0
NAND4X1
--pins(7)
Y
use :  
dir : o
shape : 
(1634,616):(1730,1584) : 0
(1604,340):(1634,1584) : 0
(1448,340):(1604,726) : 0
(1516,1412):(1604,1584) : 0
(1364,1474):(1516,1584) : 0
(1178,1474):(1364,1636) : 0
(622,1474):(1178,1584) : 0
(436,1474):(622,1636) : 0
D
use : 
dir : i
shape : 
(284,1110):(420,1272) : 0
(158,878):(284,1272) : 0
(118,878):(158,988) : 0
C
use :  
dir : i
shape : 
(670,1110):(810,1272) : 0
(546,878):(670,1272) : 0
(478,878):(546,988) : 0
B
use :  
dir : i
shape : 
(1042,1146):(1364,1324) : 0
A
use :  
dir : i
shape : 
(1290,838):(1476,1000) : 0
(838,878):(1290,988) : 0
VSS
use : g
dir : b
shape : 
(292,-160):(1800,160) : 0
(106,-160):(292,494) : 0
(0,-160):(106,160) : 0
VDD
use : p
dir : b
shape : 
(1702,2240):(1800,2560) : 0
(1516,2156):(1702,2560) : 0
(1134,2240):(1516,2560) : 0
(950,2156):(1134,2560) : 0
(284,2240):(950,2560) : 0
(98,2156):(284,2560) : 0
(0,2240):(98,2560) : 0
NAND3BXL
--pins(6)
Y
use :  
dir : o
shape : 
(1598,316):(1724,2084) : 0
(1484,316):(1598,426) : 0
(1558,1400):(1598,2084) : 0
(1516,1400):(1558,1708) : 0
(1506,1974):(1558,2084) : 0
(1004,1598):(1516,1708) : 0
(818,1572):(1004,1734) : 0
C
use : 
dir : i
shape : 
(662,1214):(786,1438) : 0
(660,1214):(662,1534) : 0
(436,1328):(660,1534) : 0
B
use :  
dir : i
shape : 
(796,758):(1162,1000) : 0
AN
use :  
dir : i
shape : 
(76,734):(284,1000) : 0
VSS
use : g
dir : b
shape : 
(644,-160):(1800,160) : 0
(458,-160):(644,244) : 0
(0,-160):(458,160) : 0
VDD
use : p
dir : b
shape : 
(1310,2240):(1800,2560) : 0
(1124,2156):(1310,2560) : 0
(644,2240):(1124,2560) : 0
(458,2156):(644,2560) : 0
(0,2240):(458,2560) : 0
NAND3BX4
--pins(6)
Y
use :  
dir : o
shape : 
(3774,398):(3900,1510) : 0
(3692,398):(3774,614) : 0
(3560,1400):(3774,1510) : 0
(1764,398):(3692,508) : 0
(3446,1400):(3560,2066) : 0
(3350,1376):(3446,2066) : 0
(3154,1376):(3350,1620) : 0
(1954,1510):(3154,1620) : 0
(1766,1484):(1954,1646) : 0
(1700,1484):(1766,1620) : 0
(1576,334):(1764,508) : 0
(1170,1510):(1700,1620) : 0
(984,1484):(1170,1646) : 0
C
use : 
dir : i
shape : 
(2468,1830):(2656,1992) : 0
(794,1858):(2468,1966) : 0
(794,878):(972,1000) : 0
(666,878):(794,1966) : 0
B
use :  
dir : i
shape : 
(2978,1014):(3166,1214) : 0
(2468,1014):(2978,1124) : 0
(2264,1014):(2468,1266) : 0
(2078,988):(2264,1266) : 0
(2064,1134):(2078,1266) : 0
(1322,1158):(2064,1266) : 0
(1134,1154):(1322,1316) : 0
AN
use :  
dir : i
shape : 
(94,822):(280,1126) : 0
VSS
use : g
dir : b
shape : 
(2810,-160):(4000,160) : 0
(2622,-160):(2810,244) : 0
(716,-160):(2622,160) : 0
(528,-160):(716,244) : 0
(0,-160):(528,160) : 0
VDD
use : p
dir : b
shape : 
(3812,2240):(4000,2560) : 0
(3686,1810):(3812,2560) : 0
(3056,2240):(3686,2560) : 0
(2868,1810):(3056,2560) : 0
(2328,2240):(2868,2560) : 0
(2140,2156):(2328,2560) : 0
(1562,2240):(2140,2560) : 0
(1374,2156):(1562,2560) : 0
(724,2240):(1374,2560) : 0
(538,2156):(724,2560) : 0
(0,2240):(538,2560) : 0
NAND3BX2
--pins(6)
Y
use :  
dir : o
shape : 
(1302,1378):(1482,1540) : 0
(1134,328):(1316,490) : 0
(1286,1378):(1302,1534) : 0
(814,1400):(1286,1534) : 0
(588,354):(1134,464) : 0
(746,1378):(814,1534) : 0
(588,1378):(746,1540) : 0
(564,354):(588,1540) : 0
(466,354):(564,1534) : 0
C
use : 
dir : i
shape : 
(2066,924):(2094,1086) : 0
(1944,924):(2066,1762) : 0
(1914,924):(1944,1086) : 0
(344,1652):(1944,1762) : 0
(222,878):(344,1762) : 0
(164,878):(222,1146) : 0
(114,878):(164,988) : 0
B
use : 
dir : i
shape : 
(1676,1014):(1740,1176) : 0
(1474,866):(1676,1208) : 0
(890,1098):(1474,1208) : 0
(710,1028):(890,1208) : 0
AN
use : #
dir : i
shape : 
(2716,934):(2726,1188) : 0
(2534,866):(2716,1188) : 0
(2524,934):(2534,1188) : 0
VSS
use : g
dir : b
shape : 
(2322,-160):(2800,160) : 0
(2290,-160):(2322,244) : 0
(2110,-160):(2290,494) : 0
(308,-160):(2110,160) : 0
(128,-160):(308,494) : 0
(0,-160):(128,160) : 0
VDD
use : p
dir : b
shape : 
(2296,2240):(2800,2560) : 0
(2116,1904):(2296,2560) : 0
(1122,2240):(2116,2560) : 0
(942,1904):(1122,2560) : 0
(384,2240):(942,2560) : 0
(204,1904):(384,2560) : 0
(0,2240):(204,2560) : 0
NAND3BX1
--pins(6)
Y
use :  
dir : o
shape : 
(1598,316):(1724,2084) : 0
(1484,316):(1598,426) : 0
(1558,1666):(1598,2084) : 0
(1004,1666):(1558,1776) : 0
(1506,1974):(1558,2084) : 0
(818,1666):(1004,1828) : 0
C
use : 
dir : i
shape : 
(660,1186):(786,1522) : 0
(478,1330):(660,1522) : 0
B
use :  
dir : i
shape : 
(796,828):(1134,1000) : 0
AN
use :  
dir : i
shape : 
(76,734):(284,1000) : 0
VSS
use : g
dir : b
shape : 
(610,-160):(1800,160) : 0
(426,-160):(610,244) : 0
(0,-160):(426,160) : 0
VDD
use : p
dir : b
shape : 
(1310,2240):(1800,2560) : 0
(1124,2156):(1310,2560) : 0
(644,2240):(1124,2560) : 0
(458,2156):(644,2560) : 0
(0,2240):(458,2560) : 0
NAND3XL
--pins(6)
Y
use :  
dir : o
shape : 
(1182,502):(1304,1564) : 0
(1124,502):(1182,664) : 0
(1124,1362):(1182,1564) : 0
(556,1454):(1124,1564) : 0
(376,1428):(556,1590) : 0
C
use : 
dir : i
shape : 
(74,974):(276,1266) : 0
B
use :  
dir : i
shape : 
(464,866):(698,1234) : 0
A
use :  
dir : i
shape : 
(1000,1072):(1058,1234) : 0
(878,612):(1000,1234) : 0
(814,612):(878,722) : 0
VSS
use : g
dir : b
shape : 
(276,-160):(1400,160) : 0
(96,-160):(276,244) : 0
(0,-160):(96,160) : 0
VDD
use : p
dir : b
shape : 
(912,2240):(1400,2560) : 0
(238,2156):(912,2560) : 0
(0,2240):(238,2560) : 0
NAND3X4
--pins(6)
Y
use :  
dir : o
shape : 
(3414,316):(3426,702) : 0
(3290,316):(3414,1488) : 0
(3240,316):(3290,702) : 0
(3020,1378):(3290,1488) : 0
(3120,316):(3240,496) : 0
(1352,386):(3120,496) : 0
(2834,1378):(3020,1540) : 0
(632,1378):(1540,1540) : 0
(644,334):(1352,496) : 0
(632,334):(644,1000) : 0
(448,334):(632,1540) : 0
(436,334):(448,1000) : 0
C
use : 
dir : i
shape : 
(2196,1054):(2226,1216) : 0
(2070,1054):(2196,1760) : 0
(2040,1054):(2070,1216) : 0
(310,1650):(2070,1760) : 0
(186,878):(310,1760) : 0
(118,878):(186,1146) : 0
B
use :  
dir : i
shape : 
(2730,988):(2790,1180) : 0
(2604,836):(2730,1180) : 0
(1854,836):(2604,946) : 0
(1670,834):(1854,996) : 0
(1642,836):(1670,996) : 0
(1516,836):(1642,1202) : 0
(954,1092):(1516,1202) : 0
(770,1028):(954,1202) : 0
A
use :  
dir : i
shape : 
(3092,852):(3158,1180) : 0
(2972,604):(3092,1180) : 0
(2968,604):(2972,998) : 0
(1352,604):(2968,714) : 0
(1228,604):(1352,984) : 0
(1168,822):(1228,984) : 0
VSS
use : g
dir : b
shape : 
(2390,-160):(3600,160) : 0
(2204,-160):(2390,244) : 0
(310,-160):(2204,160) : 0
(126,-160):(310,494) : 0
(0,-160):(126,160) : 0
VDD
use : p
dir : b
shape : 
(3390,2240):(3600,2560) : 0
(3204,1904):(3390,2560) : 0
(2648,2240):(3204,2560) : 0
(2462,1904):(2648,2560) : 0
(1912,2240):(2462,2560) : 0
(1726,1904):(1912,2560) : 0
(1154,2240):(1726,2560) : 0
(968,1904):(1154,2560) : 0
(396,2240):(968,2560) : 0
(210,1904):(396,2560) : 0
(0,2240):(210,2560) : 0
NAND3X2
--pins(6)
Y
use :  
dir : o
shape : 
(1382,1378):(1572,1540) : 0
(1204,328):(1396,490) : 0
(1364,1378):(1382,1522) : 0
(1036,1412):(1364,1522) : 0
(624,380):(1204,490) : 0
(864,1400):(1036,1540) : 0
(624,1378):(864,1540) : 0
(600,380):(624,1540) : 0
(496,380):(600,1522) : 0
C
use : 
dir : i
shape : 
(2192,1146):(2222,1412) : 0
(2062,1146):(2192,1762) : 0
(2032,1146):(2062,1412) : 0
(366,1652):(2062,1762) : 0
(334,920):(366,1762) : 0
(236,878):(334,1762) : 0
(174,878):(236,1146) : 0
(120,878):(174,988) : 0
B
use :  
dir : i
shape : 
(1814,986):(1846,1176) : 0
(1736,866):(1814,1176) : 0
(1564,866):(1736,1208) : 0
(946,1098):(1564,1208) : 0
(754,1028):(946,1208) : 0
A
use :  
dir : i
shape : 
(1204,600):(1396,980) : 0
VSS
use : g
dir : b
shape : 
(2464,-160):(2600,160) : 0
(2274,-160):(2464,244) : 0
(326,-160):(2274,160) : 0
(136,-160):(326,244) : 0
(0,-160):(136,160) : 0
VDD
use : p
dir : b
shape : 
(1190,2240):(2600,2560) : 0
(998,1904):(1190,2560) : 0
(408,2240):(998,2560) : 0
(216,1904):(408,2560) : 0
(0,2240):(216,2560) : 0
NAND3X1
--pins(6)
Y
use :  
dir : o
shape : 
(1304,1390):(1310,1624) : 0
(1182,334):(1304,1624) : 0
(1124,334):(1182,614) : 0
(1162,1390):(1182,1624) : 0
(1124,1462):(1162,1624) : 0
(586,1488):(1124,1598) : 0
(406,1462):(586,1624) : 0
C
use : 
dir : i
shape : 
(100,850):(282,1180) : 0
B
use :  
dir : i
shape : 
(464,1088):(698,1352) : 0
A
use :  
dir : i
shape : 
(1000,1002):(1058,1164) : 0
(878,612):(1000,1164) : 0
(814,612):(878,722) : 0
VSS
use : g
dir : b
shape : 
(308,-160):(1400,160) : 0
(128,-160):(308,244) : 0
(0,-160):(128,160) : 0
VDD
use : p
dir : b
shape : 
(966,2240):(1400,2560) : 0
(96,2156):(966,2560) : 0
(0,2240):(96,2560) : 0
NAND2BXL
--pins(5)
Y
use :  
dir : o
shape : 
(1294,612):(1324,1690) : 0
(1202,490):(1294,1690) : 0
(1114,490):(1202,722) : 0
(976,1580):(1202,1690) : 0
(814,612):(1114,722) : 0
(796,1554):(976,1716) : 0
B
use : 
dir : i
shape : 
(754,920):(782,1088) : 0
(464,878):(754,1088) : 0
(424,920):(464,1088) : 0
AN
use :  
dir : i
shape : 
(112,1802):(392,2066) : 0
VSS
use : g
dir : b
shape : 
(594,-160):(1400,160) : 0
(414,-160):(594,244) : 0
(0,-160):(414,160) : 0
VDD
use : p
dir : b
shape : 
(1272,2240):(1400,2560) : 0
(754,2156):(1272,2560) : 0
(0,2240):(754,2560) : 0
NAND2BX4
--pins(5)
Y
use :  
dir : o
shape : 
(2716,490):(2726,1266) : 0
(2534,490):(2716,1596) : 0
(2524,490):(2534,1266) : 0
(792,1434):(2534,1596) : 0
(1346,654):(2524,798) : 0
(1166,566):(1346,798) : 0
B
use : 
dir : i
shape : 
(1636,1136):(1970,1324) : 0
(960,1214):(1636,1324) : 0
(848,1146):(960,1324) : 0
(668,1136):(848,1324) : 0
AN
use :  
dir : i
shape : 
(90,962):(270,1266) : 0
VSS
use : g
dir : b
shape : 
(2026,-160):(2800,160) : 0
(1846,-160):(2026,508) : 0
(678,-160):(1846,160) : 0
(498,-160):(678,244) : 0
(0,-160):(498,160) : 0
VDD
use : p
dir : b
shape : 
(2672,2240):(2800,2560) : 0
(2492,1742):(2672,2560) : 0
(1992,2240):(2492,2560) : 0
(1810,1742):(1992,2560) : 0
(1312,2240):(1810,2560) : 0
(1132,1742):(1312,2560) : 0
(634,2240):(1132,2560) : 0
(454,1766):(634,2560) : 0
(0,2240):(454,2560) : 0
NAND2BX2
--pins(5)
Y
use :  
dir : o
shape : 
(2006,804):(2134,1540) : 0
(1756,804):(2006,914) : 0
(1788,1400):(2006,1540) : 0
(1600,1380):(1788,1542) : 0
(1752,722):(1756,914) : 0
(1624,634):(1752,914) : 0
(1388,634):(1624,742) : 0
(1544,1400):(1600,1540) : 0
(1220,1430):(1544,1540) : 0
(1200,580):(1388,742) : 0
(1078,1404):(1220,1540) : 0
(888,1404):(1078,1566) : 0
B
use : 
dir : i
shape : 
(1706,1098):(1878,1272) : 0
(934,1146):(1706,1254) : 0
(744,1120):(934,1280) : 0
AN
use :  
dir : i
shape : 
(94,904):(284,1254) : 0
VSS
use : g
dir : b
shape : 
(2100,-160):(2200,160) : 0
(1912,-160):(2100,556) : 0
(656,-160):(1912,160) : 0
(466,-160):(656,244) : 0
(0,-160):(466,160) : 0
VDD
use : p
dir : b
shape : 
(2100,2240):(2200,2560) : 0
(706,2156):(2100,2560) : 0
(0,2240):(706,2560) : 0
NAND2BX1
--pins(5)
Y
use :  
dir : o
shape : 
(1172,578):(1294,1616) : 0
(1114,578):(1172,740) : 0
(796,1508):(1172,1616) : 0
(934,600):(1114,734) : 0
(814,612):(934,722) : 0
B
use : 
dir : i
shape : 
(754,922):(782,1090) : 0
(464,878):(754,1090) : 0
(424,922):(464,1090) : 0
AN
use :  
dir : i
shape : 
(112,1802):(392,2066) : 0
VSS
use : g
dir : b
shape : 
(594,-160):(1400,160) : 0
(414,-160):(594,244) : 0
(0,-160):(414,160) : 0
VDD
use : p
dir : b
shape : 
(1272,2240):(1400,2560) : 0
(754,2156):(1272,2560) : 0
(0,2240):(754,2560) : 0
NAND2XL
--pins(5)
Y
use :  
dir : o
shape : 
(1090,588):(1104,1540) : 0
(1070,562):(1090,1540) : 0
(964,562):(1070,1596) : 0
(884,562):(964,724) : 0
(904,1390):(964,1596) : 0
(710,1486):(904,1596) : 0
(504,1486):(710,1648) : 0
B
use : 
dir : i
shape : 
(84,1000):(316,1290) : 0
A
use :  
dir : i
shape : 
(758,988):(824,1248) : 0
(618,878):(758,1248) : 0
(530,878):(618,988) : 0
VSS
use : g
dir : b
shape : 
(316,-160):(1200,160) : 0
(110,-160):(316,244) : 0
(0,-160):(110,160) : 0
VDD
use : p
dir : b
shape : 
(642,2240):(1200,2560) : 0
(296,2156):(642,2560) : 0
(0,2240):(296,2560) : 0
NAND2X4
--pins(5)
Y
use :  
dir : o
shape : 
(2498,490):(2522,1266) : 0
(2308,490):(2498,1596) : 0
(1058,614):(2308,758) : 0
(462,1434):(2308,1596) : 0
(866,566):(1058,758) : 0
B
use : 
dir : i
shape : 
(1688,1152):(1720,1314) : 0
(1528,1152):(1688,1324) : 0
(622,1214):(1528,1324) : 0
(368,1146):(622,1324) : 0
(338,1146):(368,1308) : 0
A
use :  
dir : i
shape : 
(2048,934):(2178,1304) : 0
(1936,934):(2048,1146) : 0
(1390,934):(1936,1042) : 0
(1210,878):(1390,1042) : 0
(1052,934):(1210,1042) : 0
(892,934):(1052,1104) : 0
(862,942):(892,1104) : 0
VSS
use : g
dir : b
shape : 
(1778,-160):(2600,160) : 0
(1588,-160):(1778,474) : 0
(348,-160):(1588,160) : 0
(158,-160):(348,244) : 0
(0,-160):(158,160) : 0
VDD
use : p
dir : b
shape : 
(2454,2240):(2600,2560) : 0
(2262,1742):(2454,2560) : 0
(1734,2240):(2262,2560) : 0
(1542,1742):(1734,2560) : 0
(1012,2240):(1542,2560) : 0
(822,1742):(1012,2560) : 0
(292,2240):(822,2560) : 0
(102,1742):(292,2560) : 0
(0,2240):(102,2560) : 0
NAND2X2
--pins(5)
Y
use :  
dir : o
shape : 
(1590,804):(1716,1540) : 0
(1360,804):(1590,914) : 0
(1558,1408):(1590,1540) : 0
(502,1408):(1558,1516) : 0
(1236,498):(1360,914) : 0
(1198,498):(1236,612) : 0
(1004,498):(1198,608) : 0
(818,446):(1004,608) : 0
B
use : 
dir : i
shape : 
(1336,1116):(1462,1290) : 0
(602,1154):(1336,1264) : 0
(400,1146):(602,1264) : 0
(370,1146):(400,1254) : 0
A
use :  
dir : i
shape : 
(796,800):(1102,1040) : 0
VSS
use : g
dir : b
shape : 
(1702,-160):(1800,160) : 0
(1516,-160):(1702,578) : 0
(284,-160):(1516,160) : 0
(98,-160):(284,244) : 0
(0,-160):(98,160) : 0
VDD
use : p
dir : b
shape : 
(1702,2240):(1800,2560) : 0
(420,2156):(1702,2560) : 0
(0,2240):(420,2560) : 0
NAND2X1
--pins(5)
Y
use :  
dir : o
shape : 
(1090,600):(1128,1486) : 0
(988,564):(1090,1486) : 0
(884,564):(988,734) : 0
(704,1376):(988,1486) : 0
(496,1376):(704,1538) : 0
B
use : 
dir : i
shape : 
(84,876):(316,1196) : 0
A
use :  
dir : i
shape : 
(484,1060):(842,1266) : 0
VSS
use : g
dir : b
shape : 
(316,-160):(1200,160) : 0
(110,-160):(316,656) : 0
(0,-160):(110,160) : 0
VDD
use : p
dir : b
shape : 
(718,2240):(1200,2560) : 0
(110,2156):(718,2560) : 0
(0,2240):(110,2560) : 0
MXI4X4
--pins(9)
Y
use :  
dir : o
shape : 
(8202,470):(8374,1808) : 0
(8170,366):(8202,2030) : 0
(8022,366):(8170,752) : 0
(8022,1422):(8170,2030) : 0
S1
use : 
dir : i
shape : 
(6410,1100):(6710,1280) : 0
S0
use :  
dir : i
shape : 
(2186,866):(2410,1134) : 0
D
use :  
dir : i
shape : 
(3000,866):(3094,1000) : 0
(2798,866):(3000,1092) : 0
C
use :  
dir : i
shape : 
(4582,600):(4824,734) : 0
(4462,600):(4582,1122) : 0
(4458,612):(4462,1122) : 0
(4406,948):(4458,1122) : 0
B
use :  
dir : i
shape : 
(2038,938):(2050,1092) : 0
(1834,604):(2038,1092) : 0
A
use :  
dir : i
shape : 
(74,1052):(416,1266) : 0
VSS
use : g
dir : b
shape : 
(8608,-160):(8800,160) : 0
(8426,-160):(8608,244) : 0
(7798,-160):(8426,160) : 0
(7616,-160):(7798,244) : 0
(7018,-160):(7616,160) : 0
(6838,-160):(7018,244) : 0
(4718,-160):(6838,160) : 0
(4536,-160):(4718,434) : 0
(2930,-160):(4536,160) : 0
(2750,-160):(2930,460) : 0
(2118,-160):(2750,160) : 0
(1936,-160):(2118,440) : 0
(304,-160):(1936,160) : 0
(122,-160):(304,578) : 0
(0,-160):(122,160) : 0
VDD
use : p
dir : b
shape : 
(8608,2240):(8800,2560) : 0
(8426,2156):(8608,2560) : 0
(7798,2240):(8426,2560) : 0
(7616,2156):(7798,2560) : 0
(6922,2240):(7616,2560) : 0
(6742,2156):(6922,2560) : 0
(4718,2240):(6742,2560) : 0
(4536,2156):(4718,2560) : 0
(2926,2240):(4536,2560) : 0
(2744,1996):(2926,2560) : 0
(2118,2240):(2744,2560) : 0
(1936,1996):(2118,2560) : 0
(304,2240):(1936,2560) : 0
(122,1732):(304,2560) : 0
(0,2240):(122,2560) : 0
MXI4X2
--pins(9)
Y
use :  
dir : o
shape : 
(8174,366):(8296,2014) : 0
(8104,366):(8174,752) : 0
(8164,1254):(8174,2014) : 0
(8098,1330):(8164,2014) : 0
(7774,1330):(8098,1534) : 0
S1
use : 
dir : i
shape : 
(6374,866):(6742,1048) : 0
S0
use :  
dir : i
shape : 
(2106,866):(2376,1134) : 0
D
use :  
dir : i
shape : 
(2874,604):(3096,1066) : 0
C
use :  
dir : i
shape : 
(4584,600):(4826,734) : 0
(4466,600):(4584,1122) : 0
(4462,612):(4466,1122) : 0
(4410,948):(4462,1122) : 0
B
use :  
dir : i
shape : 
(1938,612):(1986,722) : 0
(1816,612):(1938,1054) : 0
(1724,900):(1816,1054) : 0
A
use :  
dir : i
shape : 
(74,1052):(418,1266) : 0
VSS
use : g
dir : b
shape : 
(7848,-160):(8400,160) : 0
(7668,-160):(7848,244) : 0
(6936,-160):(7668,160) : 0
(6756,-160):(6936,244) : 0
(4720,-160):(6756,160) : 0
(4540,-160):(4720,434) : 0
(3044,-160):(4540,160) : 0
(2864,-160):(3044,434) : 0
(2084,-160):(2864,160) : 0
(1904,-160):(2084,440) : 0
(302,-160):(1904,160) : 0
(122,-160):(302,658) : 0
(0,-160):(122,160) : 0
VDD
use : p
dir : b
shape : 
(7800,2240):(8400,2560) : 0
(7620,2156):(7800,2560) : 0
(6868,2240):(7620,2560) : 0
(6688,2156):(6868,2560) : 0
(4720,2240):(6688,2560) : 0
(4540,2156):(4720,2560) : 0
(2938,2240):(4540,2560) : 0
(2758,1908):(2938,2560) : 0
(2084,2240):(2758,2560) : 0
(1904,1908):(2084,2560) : 0
(302,2240):(1904,2560) : 0
(122,1490):(302,2560) : 0
(0,2240):(122,2560) : 0
MXI2X4
--pins(6)
Y
use :  
dir : o
shape : 
(3036,342):(3208,524) : 0
(2310,1708):(3054,1816) : 0
(2430,342):(3036,452) : 0
(2424,342):(2430,510) : 0
(2310,334):(2424,1000) : 0
(2218,334):(2310,1816) : 0
(1656,342):(2218,452) : 0
(2186,878):(2218,1816) : 0
(2026,1666):(2186,1816) : 0
(1388,1708):(2026,1816) : 0
(1472,342):(1656,504) : 0
S0
use : 
dir : i
shape : 
(3204,1908):(3388,2070) : 0
(2932,1934):(3204,2070) : 0
(1252,1960):(2932,2070) : 0
(1128,1886):(1252,2070) : 0
B
use : 
dir : i
shape : 
(4004,1028):(4378,1266) : 0
A
use : �
dir : i
shape : 
(598,1052):(812,1214) : 0
(474,1052):(598,1254) : 0
(304,1052):(474,1214) : 0
VSS
use : g
dir : b
shape : 
(4902,-160):(5000,160) : 0
(4718,-160):(4902,470) : 0
(4156,-160):(4718,160) : 0
(3972,-160):(4156,244) : 0
(998,-160):(3972,160) : 0
(814,-160):(998,470) : 0
(292,-160):(814,160) : 0
(108,-160):(292,480) : 0
(0,-160):(108,160) : 0
VDD
use : p
dir : b
shape : 
(4902,2240):(5000,2560) : 0
(4718,1958):(4902,2560) : 0
(4142,2240):(4718,2560) : 0
(3958,1792):(4142,2560) : 0
(966,2240):(3958,2560) : 0
(842,1958):(966,2560) : 0
(292,2240):(842,2560) : 0
(108,1964):(292,2560) : 0
(0,2240):(108,2560) : 0
MXI2X2
--pins(6)
Y
use :  
dir : o
shape : 
(1766,586):(1888,1776) : 0
(1676,1666):(1766,1776) : 0
(1432,1666):(1676,2010) : 0
S0
use : 
dir : i
shape : 
(358,1312):(626,1534) : 0
B
use :  
dir : i
shape : 
(774,1012):(986,1266) : 0
A
use :  
dir : i
shape : 
(2504,866):(2726,1152) : 0
VSS
use : g
dir : b
shape : 
(2704,-160):(2800,160) : 0
(2524,-160):(2704,244) : 0
(918,-160):(2524,160) : 0
(738,-160):(918,522) : 0
(0,-160):(738,160) : 0
VDD
use : p
dir : b
shape : 
(2704,2240):(2800,2560) : 0
(2524,1514):(2704,2560) : 0
(754,2240):(2524,2560) : 0
(572,1706):(754,2560) : 0
(0,2240):(572,2560) : 0
MXI2X1
--pins(6)
Y
use :  
dir : o
shape : 
(1658,1146):(1736,1610) : 0
(1658,562):(1688,724) : 0
(1528,562):(1658,1610) : 0
(1496,562):(1528,724) : 0
(1496,1448):(1528,1610) : 0
S0
use : 
dir : i
shape : 
(396,1048):(664,1266) : 0
B
use :  
dir : i
shape : 
(822,866):(1058,1110) : 0
A
use :  
dir : i
shape : 
(2256,866):(2522,1086) : 0
VSS
use : g
dir : b
shape : 
(2494,-160):(2600,160) : 0
(2302,-160):(2494,244) : 0
(822,-160):(2302,160) : 0
(630,-160):(822,694) : 0
(0,-160):(630,160) : 0
VDD
use : p
dir : b
shape : 
(2502,2240):(2600,2560) : 0
(2304,2128):(2502,2560) : 0
(800,2240):(2304,2560) : 0
(608,1908):(800,2560) : 0
(0,2240):(608,2560) : 0
MX4X4
--pins(9)
Y
use :  
dir : o
shape : 
(7774,640):(7976,1800) : 0
(7730,640):(7774,848) : 0
(7730,1314):(7774,1800) : 0
S1
use : 
dir : i
shape : 
(6860,1158):(7026,1320) : 0
(6738,1158):(6860,1788) : 0
(5876,1678):(6738,1788) : 0
(5674,1678):(5876,1838) : 0
S0
use :  
dir : i
shape : 
(4048,1902):(4170,2066) : 0
(1514,1902):(4048,2012) : 0
(1286,1902):(1514,2028) : 0
(1260,1902):(1286,2054) : 0
(1236,1920):(1260,2054) : 0
(1056,1920):(1236,2080) : 0
D
use :  
dir : i
shape : 
(2214,1122):(2336,1254) : 0
(2020,1122):(2214,1230) : 0
(1898,1048):(2020,1230) : 0
C
use :  
dir : i
shape : 
(222,866):(404,1100) : 0
(74,866):(222,1098) : 0
B
use :  
dir : i
shape : 
(3160,866):(3426,1080) : 0
A
use :  
dir : i
shape : 
(4906,1050):(5176,1266) : 0
VSS
use : g
dir : b
shape : 
(8256,-160):(8400,160) : 0
(8076,-160):(8256,484) : 0
(7556,-160):(8076,160) : 0
(7376,-160):(7556,448) : 0
(5216,-160):(7376,160) : 0
(5036,-160):(5216,244) : 0
(3218,-160):(5036,160) : 0
(3038,-160):(3218,244) : 0
(2290,-160):(3038,160) : 0
(2110,-160):(2290,244) : 0
(276,-160):(2110,160) : 0
(96,-160):(276,728) : 0
(0,-160):(96,160) : 0
VDD
use : p
dir : b
shape : 
(8256,2240):(8400,2560) : 0
(8076,1964):(8256,2560) : 0
(7556,2240):(8076,2560) : 0
(7376,1964):(7556,2560) : 0
(5212,2240):(7376,2560) : 0
(5032,2156):(5212,2560) : 0
(3218,2240):(5032,2560) : 0
(3038,2156):(3218,2560) : 0
(2224,2240):(3038,2560) : 0
(2044,2156):(2224,2560) : 0
(276,2240):(2044,2560) : 0
(96,1514):(276,2560) : 0
(0,2240):(96,2560) : 0
MX4X2
--pins(9)
Y
use :  
dir : o
shape : 
(7812,1412):(7886,1522) : 0
(7692,360):(7812,2012) : 0
(7634,360):(7692,746) : 0
(7634,1402):(7692,2012) : 0
S1
use : 
dir : i
shape : 
(6816,1158):(6982,1320) : 0
(6696,1158):(6816,1788) : 0
(5840,1678):(6696,1788) : 0
(5638,1678):(5840,1838) : 0
S0
use :  
dir : i
shape : 
(4024,1902):(4144,2066) : 0
(1504,1902):(4024,2012) : 0
(1278,1902):(1504,2028) : 0
(1252,1902):(1278,2054) : 0
(1228,1920):(1252,2054) : 0
(1048,1920):(1228,2080) : 0
D
use :  
dir : i
shape : 
(2200,1122):(2322,1254) : 0
(2008,1122):(2200,1230) : 0
(1886,1048):(2008,1230) : 0
C
use :  
dir : i
shape : 
(222,866):(400,1100) : 0
(74,866):(222,1098) : 0
B
use :  
dir : i
shape : 
(3140,866):(3404,1080) : 0
A
use :  
dir : i
shape : 
(4874,1050):(5144,1266) : 0
VSS
use : g
dir : b
shape : 
(7402,-160):(8000,160) : 0
(7222,-160):(7402,420) : 0
(5184,-160):(7222,160) : 0
(5004,-160):(5184,244) : 0
(3198,-160):(5004,160) : 0
(3020,-160):(3198,244) : 0
(2276,-160):(3020,160) : 0
(2098,-160):(2276,244) : 0
(274,-160):(2098,160) : 0
(94,-160):(274,728) : 0
(0,-160):(94,160) : 0
VDD
use : p
dir : b
shape : 
(7402,2240):(8000,2560) : 0
(7222,1754):(7402,2560) : 0
(5180,2240):(7222,2560) : 0
(5002,2156):(5180,2560) : 0
(3198,2240):(5002,2560) : 0
(3020,2156):(3198,2560) : 0
(2210,2240):(3020,2560) : 0
(2032,2156):(2210,2560) : 0
(274,2240):(2032,2560) : 0
(94,1514):(274,2560) : 0
(0,2240):(94,2560) : 0
MX2X4
--pins(6)
Y
use :  
dir : o
shape : 
(2956,334):(3164,1596) : 0
(2848,1414):(2956,1596) : 0
S0
use : 
dir : i
shape : 
(532,1400):(1004,1534) : 0
(340,1354):(532,1534) : 0
B
use :  
dir : i
shape : 
(470,842):(826,1024) : 0
(436,866):(470,1024) : 0
A
use :  
dir : i
shape : 
(2236,866):(2522,1066) : 0
VSS
use : g
dir : b
shape : 
(3496,-160):(3600,160) : 0
(3310,-160):(3496,422) : 0
(2744,-160):(3310,160) : 0
(2558,-160):(2744,422) : 0
(796,-160):(2558,160) : 0
(610,-160):(796,704) : 0
(0,-160):(610,160) : 0
VDD
use : p
dir : b
shape : 
(3490,2240):(3600,2560) : 0
(3306,2156):(3490,2560) : 0
(2640,2240):(3306,2560) : 0
(2454,1972):(2640,2560) : 0
(710,2240):(2454,2560) : 0
(524,1710):(710,2560) : 0
(0,2240):(524,2560) : 0
MX2X2
--pins(6)
Y
use :  
dir : o
shape : 
(2988,388):(3112,1954) : 0
(2960,388):(2988,878) : 0
(2892,1400):(2988,1954) : 0
(2922,388):(2960,790) : 0
S0
use : 
dir : i
shape : 
(604,1412):(950,1522) : 0
(450,1412):(604,1590) : 0
(420,1428):(450,1590) : 0
B
use :  
dir : i
shape : 
(430,1052):(774,1266) : 0
A
use :  
dir : i
shape : 
(2570,612):(2728,722) : 0
(2444,612):(2570,734) : 0
(2320,612):(2444,1150) : 0
VSS
use : g
dir : b
shape : 
(2672,-160):(3200,160) : 0
(2488,-160):(2672,446) : 0
(814,-160):(2488,160) : 0
(630,-160):(814,592) : 0
(0,-160):(630,160) : 0
VDD
use : p
dir : b
shape : 
(2646,2240):(3200,2560) : 0
(2462,2156):(2646,2560) : 0
(814,2240):(2462,2560) : 0
(630,1780):(814,2560) : 0
(0,2240):(630,2560) : 0
MX2X1
--pins(6)
Y
use :  
dir : o
shape : 
(2604,536):(2726,1892) : 0
(2500,536):(2604,758) : 0
(2396,1508):(2604,1892) : 0
(2496,536):(2500,722) : 0
S0
use : 
dir : i
shape : 
(74,1888):(376,2066) : 0
B
use :  
dir : i
shape : 
(774,1376):(976,1534) : 0
(584,1270):(774,1534) : 0
A
use :  
dir : i
shape : 
(2000,866):(2376,1054) : 0
VSS
use : g
dir : b
shape : 
(2278,-160):(2800,160) : 0
(2098,-160):(2278,244) : 0
(698,-160):(2098,160) : 0
(698,582):(702,684) : 0
(528,-160):(698,684) : 0
(0,-160):(528,160) : 0
(522,582):(528,684) : 0
VDD
use : p
dir : b
shape : 
(2280,2240):(2800,2560) : 0
(2100,2156):(2280,2560) : 0
(678,2240):(2100,2560) : 0
(498,1704):(678,2560) : 0
(0,2240):(498,2560) : 0
INVXL
--pins(4)
Y
use :  
dir : o
shape : 
(624,1134):(716,1536) : 0
(624,642):(678,878) : 0
(484,642):(624,1536) : 0
(472,642):(484,878) : 0
A
use : 
dir : i
shape : 
(84,866):(316,1196) : 0
VSS
use : g
dir : b
shape : 
(600,-160):(800,160) : 0
(110,-160):(600,244) : 0
(0,-160):(110,160) : 0
VDD
use : p
dir : b
shape : 
(516,2240):(800,2560) : 0
(516,1850):(658,1950) : 0
(310,1850):(516,2560) : 0
(166,1850):(310,1950) : 0
(0,2240):(310,2560) : 0
INVX8
--pins(4)
Y
use :  
dir : o
shape : 
(1756,838):(2080,1534) : 0
(1714,722):(1756,1534) : 0
(1622,722):(1714,1560) : 0
(1220,614):(1622,1624) : 0
(1178,614):(1220,866) : 0
(434,1396):(1220,1624) : 0
(434,614):(1178,842) : 0
A
use : 
dir : i
shape : 
(300,974):(752,1266) : 0
VSS
use : g
dir : b
shape : 
(2086,-160):(2200,160) : 0
(1636,-160):(2086,244) : 0
(1066,-160):(1636,160) : 0
(878,-160):(1066,428) : 0
(312,-160):(878,160) : 0
(122,-160):(312,244) : 0
(0,-160):(122,160) : 0
VDD
use : p
dir : b
shape : 
(2100,2240):(2200,2560) : 0
(1844,2156):(2100,2560) : 0
(1656,1834):(1844,2560) : 0
(1064,2240):(1656,2560) : 0
(876,1834):(1064,2560) : 0
(288,2240):(876,2560) : 0
(100,1834):(288,2560) : 0
(0,2240):(100,2560) : 0
INVX4
--pins(4)
Y
use :  
dir : o
shape : 
(502,388):(682,2020) : 0
(424,866):(502,1534) : 0
A
use : 
dir : i
shape : 
(74,892):(276,1266) : 0
VSS
use : g
dir : b
shape : 
(1084,-160):(1400,160) : 0
(904,-160):(1084,744) : 0
(276,-160):(904,160) : 0
(96,-160):(276,744) : 0
(0,-160):(96,160) : 0
VDD
use : p
dir : b
shape : 
(1084,2240):(1400,2560) : 0
(904,1440):(1084,2560) : 0
(276,2240):(904,2560) : 0
(96,1440):(276,2560) : 0
(0,2240):(96,2560) : 0
INVX2
--pins(4)
Y
use :  
dir : o
shape : 
(976,366):(1116,1430) : 0
(884,366):(976,752) : 0
(930,1254):(976,1430) : 0
(654,1322):(930,1430) : 0
(448,1322):(654,1708) : 0
A
use : 
dir : i
shape : 
(300,866):(790,1148) : 0
VSS
use : g
dir : b
shape : 
(534,-160):(1200,160) : 0
(328,-160):(534,722) : 0
(0,-160):(328,160) : 0
VDD
use : p
dir : b
shape : 
(994,2240):(1200,2560) : 0
(990,2156):(994,2560) : 0
(790,2128):(990,2560) : 0
(788,2156):(790,2560) : 0
(0,2240):(788,2560) : 0
INVX20
--pins(4)
Y
use :  
dir : o
shape : 
(5672,570):(6486,1828) : 0
(5466,570):(5672,896) : 0
(5386,1424):(5672,1748) : 0
(3798,572):(5466,896) : 0
(5098,1392):(5386,1778) : 0
(4640,1424):(5098,1748) : 0
(4402,1392):(4640,1778) : 0
(3934,1424):(4402,1748) : 0
(3708,1392):(3934,1778) : 0
(3618,570):(3798,896) : 0
(3240,1424):(3708,1748) : 0
(2960,570):(3618,892) : 0
(2960,1392):(3240,1778) : 0
A
use : 
dir : i
shape : 
(422,1000):(660,1266) : 0
VSS
use : g
dir : b
shape : 
(6492,-160):(6600,160) : 0
(6314,-160):(6492,244) : 0
(5764,-160):(6314,160) : 0
(5584,-160):(5764,244) : 0
(5016,-160):(5584,160) : 0
(4836,-160):(5016,244) : 0
(4264,-160):(4836,160) : 0
(4084,-160):(4264,244) : 0
(3516,-160):(4084,160) : 0
(3336,-160):(3516,244) : 0
(2782,-160):(3336,160) : 0
(2602,-160):(2782,244) : 0
(2022,-160):(2602,160) : 0
(1842,-160):(2022,456) : 0
(1272,-160):(1842,160) : 0
(1092,-160):(1272,456) : 0
(528,-160):(1092,160) : 0
(350,-160):(528,772) : 0
(0,-160):(350,160) : 0
VDD
use : p
dir : b
shape : 
(6492,2240):(6600,2560) : 0
(6314,2156):(6492,2560) : 0
(5764,2240):(6314,2560) : 0
(5584,2156):(5764,2560) : 0
(5016,2240):(5584,2560) : 0
(4836,2156):(5016,2560) : 0
(4260,2240):(4836,2560) : 0
(4082,2156):(4260,2560) : 0
(3514,2240):(4082,2560) : 0
(3334,2156):(3514,2560) : 0
(2768,2240):(3334,2560) : 0
(2590,2156):(2768,2560) : 0
(2018,2240):(2590,2560) : 0
(1840,1964):(2018,2560) : 0
(1244,2240):(1840,2560) : 0
(1066,1978):(1244,2560) : 0
(528,2240):(1066,2560) : 0
(350,1482):(528,2560) : 0
(0,2240):(350,2560) : 0
INVX1
--pins(4)
Y
use :  
dir : o
shape : 
(646,1128):(716,1696) : 0
(506,642):(646,1696) : 0
(484,1128):(506,1696) : 0
A
use : 
dir : i
shape : 
(84,866):(346,1136) : 0
VSS
use : g
dir : b
shape : 
(316,-160):(800,160) : 0
(110,-160):(316,244) : 0
(0,-160):(110,160) : 0
VDD
use : p
dir : b
shape : 
(316,2240):(800,2560) : 0
(110,2156):(316,2560) : 0
(0,2240):(110,2560) : 0
INVX16
--pins(4)
Y
use :  
dir : o
shape : 
(5056,572):(5886,1828) : 0
(3858,572):(5056,896) : 0
(4714,1424):(5056,1748) : 0
(4474,1392):(4714,1778) : 0
(3998,1424):(4474,1748) : 0
(3768,1392):(3998,1778) : 0
(3676,570):(3858,896) : 0
(3292,1424):(3768,1748) : 0
(3008,570):(3676,892) : 0
(3008,1392):(3292,1778) : 0
A
use : 
dir : i
shape : 
(428,1000):(672,1266) : 0
VSS
use : g
dir : b
shape : 
(5856,-160):(6000,160) : 0
(5674,-160):(5856,244) : 0
(5096,-160):(5674,160) : 0
(4914,-160):(5096,244) : 0
(4332,-160):(4914,160) : 0
(4150,-160):(4332,244) : 0
(3570,-160):(4150,160) : 0
(3388,-160):(3570,244) : 0
(2826,-160):(3388,160) : 0
(2644,-160):(2826,244) : 0
(2054,-160):(2644,160) : 0
(1872,-160):(2054,456) : 0
(1292,-160):(1872,160) : 0
(1110,-160):(1292,456) : 0
(516,-160):(1110,160) : 0
(334,-160):(516,818) : 0
(0,-160):(334,160) : 0
VDD
use : p
dir : b
shape : 
(5856,2240):(6000,2560) : 0
(5674,2156):(5856,2560) : 0
(5096,2240):(5674,2560) : 0
(4914,2156):(5096,2560) : 0
(4328,2240):(4914,2560) : 0
(4148,2156):(4328,2560) : 0
(3570,2240):(4148,2560) : 0
(3388,2156):(3570,2560) : 0
(2818,2240):(3388,2560) : 0
(2636,2156):(2818,2560) : 0
(2050,2240):(2636,2560) : 0
(1868,1964):(2050,2560) : 0
(1264,2240):(1868,2560) : 0
(1082,1978):(1264,2560) : 0
(516,2240):(1082,2560) : 0
(334,1482):(516,2560) : 0
(0,2240):(334,2560) : 0
INVX12
--pins(4)
Y
use :  
dir : o
shape : 
(3654,572):(4484,1828) : 0
(2310,572):(3654,896) : 0
(3614,1252):(3654,1828) : 0
(2308,1352):(3614,1828) : 0
A
use : 
dir : i
shape : 
(278,1014):(462,1176) : 0
(238,1066):(278,1176) : 0
(116,1066):(238,1254) : 0
VSS
use : g
dir : b
shape : 
(4498,-160):(4600,160) : 0
(4316,-160):(4498,398) : 0
(3736,-160):(4316,160) : 0
(3554,-160):(3736,398) : 0
(2968,-160):(3554,160) : 0
(2786,-160):(2968,398) : 0
(1490,-160):(2786,160) : 0
(1308,-160):(1490,244) : 0
(748,-160):(1308,160) : 0
(566,-160):(748,474) : 0
(0,-160):(566,160) : 0
VDD
use : p
dir : b
shape : 
(4504,2240):(4600,2560) : 0
(4322,1978):(4504,2560) : 0
(3736,2240):(4322,2560) : 0
(3554,1978):(3736,2560) : 0
(2968,2240):(3554,2560) : 0
(2786,1978):(2968,2560) : 0
(2220,2240):(2786,2560) : 0
(2034,2130):(2220,2560) : 0
(718,2240):(2034,2560) : 0
(536,2156):(718,2560) : 0
(0,2240):(536,2560) : 0
DFFRHQX1
--pins(6)
RN
use :  
dir : i
shape : 
(6198,1386):(6620,1552) : 0
Q
use : 
dir : o
shape : 
(7278,592):(7286,1522) : 0
(7162,592):(7278,2042) : 0
(6712,592):(7162,702) : 0
(7122,1412):(7162,2042) : 0
(7096,1658):(7122,2042) : 0
(6588,348):(6712,702) : 0
(6530,348):(6588,510) : 0
D
use : 
dir : i
shape : 
(862,612):(942,722) : 0
(862,862):(864,1024) : 0
(740,612):(862,1024) : 0
(684,862):(740,1024) : 0
CK
use : c
dir : i
shape : 
(480,1146):(590,1266) : 0
(310,1034):(480,1266) : 0
VSS
use : g
dir : b
shape : 
(7096,-160):(7400,160) : 0
(6914,-160):(7096,422) : 0
(6302,-160):(6914,160) : 0
(5800,-160):(6302,244) : 0
(5192,-160):(5800,160) : 0
(5010,-160):(5192,244) : 0
(3628,-160):(5010,160) : 0
(3446,-160):(3628,508) : 0
(2146,-160):(3446,160) : 0
(1964,-160):(2146,654) : 0
(692,-160):(1964,160) : 0
(510,-160):(692,468) : 0
(0,-160):(510,160) : 0
VDD
use : p
dir : b
shape : 
(6594,2240):(7400,2560) : 0
(6412,1706):(6594,2560) : 0
(5388,2240):(6412,2560) : 0
(5166,2156):(5388,2560) : 0
(3852,2240):(5166,2560) : 0
(3630,2156):(3852,2560) : 0
(2156,2240):(3630,2560) : 0
(1976,1926):(2156,2560) : 0
(844,2240):(1976,2560) : 0
(662,1840):(844,2560) : 0
(0,2240):(662,2560) : 0
CLKINVX8
--pins(4)
Y
use :  
dir : o
shape : 
(1756,866):(2080,1534) : 0
(1714,720):(1756,1534) : 0
(1600,720):(1714,1560) : 0
(1220,588):(1600,1624) : 0
(1178,588):(1220,866) : 0
(434,1396):(1220,1624) : 0
(484,588):(1178,816) : 0
A
use : 
dir : i
shape : 
(300,974):(752,1266) : 0
VSS
use : g
dir : b
shape : 
(1114,-160):(2200,160) : 0
(926,-160):(1114,436) : 0
(312,-160):(926,160) : 0
(122,-160):(312,244) : 0
(0,-160):(122,160) : 0
VDD
use : p
dir : b
shape : 
(1844,2240):(2200,2560) : 0
(1656,1834):(1844,2560) : 0
(1064,2240):(1656,2560) : 0
(876,1834):(1064,2560) : 0
(288,2240):(876,2560) : 0
(100,1834):(288,2560) : 0
(0,2240):(100,2560) : 0
CLKINVX4
--pins(4)
Y
use :  
dir : o
shape : 
(774,614):(976,1800) : 0
(572,614):(774,796) : 0
(764,1412):(774,1800) : 0
(584,1412):(764,2002) : 0
A
use : 
dir : i
shape : 
(74,962):(504,1266) : 0
VSS
use : g
dir : b
shape : 
(1294,-160):(1400,160) : 0
(1114,-160):(1294,244) : 0
(360,-160):(1114,160) : 0
(180,-160):(360,244) : 0
(0,-160):(180,160) : 0
VDD
use : p
dir : b
shape : 
(1166,2240):(1400,2560) : 0
(986,2156):(1166,2560) : 0
(360,2240):(986,2560) : 0
(180,2156):(360,2560) : 0
(0,2240):(180,2560) : 0
CLKINVX3
--pins(4)
Y
use :  
dir : o
shape : 
(622,1252):(716,1800) : 0
(482,684):(622,1800) : 0
(446,1254):(482,1800) : 0
A
use : 
dir : i
shape : 
(84,866):(324,1162) : 0
VSS
use : g
dir : b
shape : 
(994,-160):(1200,160) : 0
(788,-160):(994,244) : 0
(0,-160):(788,160) : 0
VDD
use : p
dir : b
shape : 
(316,2240):(1200,2560) : 0
(110,2156):(316,2560) : 0
(0,2240):(110,2560) : 0
CLKINVX2
--pins(4)
Y
use :  
dir : o
shape : 
(800,572):(940,1574) : 0
(700,572):(800,734) : 0
(448,1400):(800,1574) : 0
A
use : 
dir : i
shape : 
(84,866):(658,1148) : 0
VSS
use : g
dir : b
shape : 
(440,-160):(1200,160) : 0
(234,-160):(440,704) : 0
(0,-160):(234,160) : 0
VDD
use : p
dir : b
shape : 
(878,2240):(1200,2560) : 0
(648,2122):(878,2560) : 0
(0,2240):(648,2560) : 0
CLKINVX20
--pins(4)
Y
use :  
dir : o
shape : 
(9734,1392):(10066,1778) : 0
(8908,572):(9734,1800) : 0
(4742,570):(8908,872) : 0
(8556,1424):(8908,1748) : 0
(8254,1392):(8556,1778) : 0
(7852,1424):(8254,1748) : 0
(7524,1392):(7852,1778) : 0
(6958,1424):(7524,1748) : 0
(6776,1392):(6958,1778) : 0
(6192,1424):(6776,1748) : 0
(5864,1392):(6192,1778) : 0
(5436,1424):(5864,1748) : 0
(5162,1392):(5436,1778) : 0
(4686,1424):(5162,1748) : 0
(4458,1392):(4686,1778) : 0
(3984,1424):(4458,1748) : 0
(3736,1392):(3984,1778) : 0
A
use : 
dir : i
shape : 
(382,1000):(628,1266) : 0
VSS
use : g
dir : b
shape : 
(8410,-160):(10200,160) : 0
(8228,-160):(8410,428) : 0
(7672,-160):(8228,160) : 0
(7490,-160):(7672,428) : 0
(6914,-160):(7490,160) : 0
(6734,-160):(6914,428) : 0
(6152,-160):(6734,160) : 0
(5972,-160):(6152,428) : 0
(5396,-160):(5972,160) : 0
(5214,-160):(5396,428) : 0
(4640,-160):(5214,160) : 0
(4458,-160):(4640,428) : 0
(2764,-160):(4458,160) : 0
(2582,-160):(2764,420) : 0
(1940,-160):(2582,160) : 0
(1758,-160):(1940,420) : 0
(1180,-160):(1758,160) : 0
(1000,-160):(1180,446) : 0
(0,-160):(1000,160) : 0
VDD
use : p
dir : b
shape : 
(9600,2240):(10200,2560) : 0
(9420,1992):(9600,2560) : 0
(8842,2240):(9420,2560) : 0
(8660,1992):(8842,2560) : 0
(8084,2240):(8660,2560) : 0
(7904,1992):(8084,2560) : 0
(7324,2240):(7904,2560) : 0
(7144,1992):(7324,2560) : 0
(6574,2240):(7144,2560) : 0
(6392,1992):(6574,2560) : 0
(5816,2240):(6392,2560) : 0
(5636,1966):(5816,2560) : 0
(5052,2240):(5636,2560) : 0
(4870,1966):(5052,2560) : 0
(4296,2240):(4870,2560) : 0
(4114,1966):(4296,2560) : 0
(3538,2240):(4114,2560) : 0
(3358,1970):(3538,2560) : 0
(2702,2240):(3358,2560) : 0
(2520,1964):(2702,2560) : 0
(1938,2240):(2520,2560) : 0
(1756,1964):(1938,2560) : 0
(1154,2240):(1756,2560) : 0
(972,1978):(1154,2560) : 0
(428,2240):(972,2560) : 0
(248,1482):(428,2560) : 0
(0,2240):(248,2560) : 0
CLKINVX16
--pins(4)
Y
use :  
dir : o
shape : 
(7858,572):(8686,1828) : 0
(6928,572):(7858,896) : 0
(7570,1424):(7858,1748) : 0
(7278,1392):(7570,1778) : 0
(6822,1424):(7278,1748) : 0
(6242,570):(6928,896) : 0
(6574,1392):(6822,1778) : 0
(6098,1424):(6574,1748) : 0
(4370,572):(6242,896) : 0
(5870,1392):(6098,1778) : 0
(5394,1424):(5870,1748) : 0
(5118,1392):(5394,1778) : 0
(4690,1424):(5118,1748) : 0
(4354,1392):(4690,1778) : 0
(3778,1424):(4354,1748) : 0
(3598,1392):(3778,1778) : 0
A
use : 
dir : i
shape : 
(382,1000):(630,1266) : 0
VSS
use : g
dir : b
shape : 
(7282,-160):(8800,160) : 0
(7102,-160):(7282,428) : 0
(6544,-160):(7102,160) : 0
(6362,-160):(6544,428) : 0
(5786,-160):(6362,160) : 0
(5606,-160):(5786,428) : 0
(5024,-160):(5606,160) : 0
(4842,-160):(5024,428) : 0
(4266,-160):(4842,160) : 0
(4086,-160):(4266,428) : 0
(1942,-160):(4086,160) : 0
(1760,-160):(1942,456) : 0
(1182,-160):(1760,160) : 0
(1000,-160):(1182,446) : 0
(0,-160):(1000,160) : 0
VDD
use : p
dir : b
shape : 
(8662,2240):(8800,2560) : 0
(8480,1992):(8662,2560) : 0
(7950,2240):(8480,2560) : 0
(7768,1992):(7950,2560) : 0
(7190,2240):(7768,2560) : 0
(7008,1992):(7190,2560) : 0
(6438,2240):(7008,2560) : 0
(6256,1992):(6438,2560) : 0
(5680,2240):(6256,2560) : 0
(5498,1966):(5680,2560) : 0
(4914,2240):(5498,2560) : 0
(4734,1966):(4914,2560) : 0
(4158,2240):(4734,2560) : 0
(3976,1966):(4158,2560) : 0
(3400,2240):(3976,2560) : 0
(3218,1970):(3400,2560) : 0
(2704,2240):(3218,2560) : 0
(2522,1964):(2704,2560) : 0
(1938,2240):(2522,2560) : 0
(1758,1964):(1938,2560) : 0
(1154,2240):(1758,2560) : 0
(974,1978):(1154,2560) : 0
(430,2240):(974,2560) : 0
(248,1482):(430,2560) : 0
(0,2240):(248,2560) : 0
CLKBUFXL
--pins(4)
Y
use :  
dir : o
shape : 
(1164,580):(1286,1424) : 0
(1018,580):(1164,690) : 0
(1124,1254):(1164,1424) : 0
(996,1314):(1124,1424) : 0
(838,528):(1018,690) : 0
(816,1314):(996,1476) : 0
A
use : 
dir : i
shape : 
(74,836):(430,1070) : 0
VSS
use : g
dir : b
shape : 
(594,-160):(1400,160) : 0
(414,-160):(594,244) : 0
(0,-160):(414,160) : 0
VDD
use : p
dir : b
shape : 
(646,2240):(1400,2560) : 0
(466,2156):(646,2560) : 0
(0,2240):(466,2560) : 0
CLKBUFX8
--pins(4)
Y
use :  
dir : o
shape : 
(2252,866):(2480,1534) : 0
(1606,642):(2252,1534) : 0
(1564,642):(1606,880) : 0
(1564,1250):(1606,1514) : 0
(1272,642):(1564,804) : 0
(1226,1352):(1564,1514) : 0
A
use : 
dir : i
shape : 
(622,948):(782,1110) : 0
(492,878):(622,1110) : 0
(320,948):(492,1110) : 0
VSS
use : g
dir : b
shape : 
(1824,-160):(2600,160) : 0
(1632,-160):(1824,430) : 0
(1104,-160):(1632,160) : 0
(912,-160):(1104,430) : 0
(0,-160):(912,160) : 0
VDD
use : p
dir : b
shape : 
(2498,2240):(2600,2560) : 0
(2308,1754):(2498,2560) : 0
(1778,2240):(2308,2560) : 0
(1588,1754):(1778,2560) : 0
(1036,2240):(1588,2560) : 0
(844,2156):(1036,2560) : 0
(292,2240):(844,2560) : 0
(102,1688):(292,2560) : 0
(0,2240):(102,2560) : 0
CLKBUFX4
--pins(4)
Y
use :  
dir : o
shape : 
(1282,600):(1364,1266) : 0
(1156,600):(1282,1428) : 0
(928,662):(1156,824) : 0
(1112,1320):(1156,1428) : 0
(928,1320):(1112,1480) : 0
A
use : 
dir : i
shape : 
(76,866):(442,1140) : 0
VSS
use : g
dir : b
shape : 
(1528,-160):(1800,160) : 0
(1342,-160):(1528,244) : 0
(644,-160):(1342,160) : 0
(458,-160):(644,244) : 0
(0,-160):(458,160) : 0
VDD
use : p
dir : b
shape : 
(1528,2240):(1800,2560) : 0
(1342,2156):(1528,2560) : 0
(698,2240):(1342,2560) : 0
(668,2156):(698,2560) : 0
(542,2130):(668,2560) : 0
(512,2156):(542,2560) : 0
(0,2240):(512,2560) : 0
CLKBUFX3
--pins(4)
Y
use :  
dir : o
shape : 
(938,574):(996,736) : 0
(938,866):(976,1504) : 0
(816,574):(938,1504) : 0
(796,866):(816,1504) : 0
(774,866):(796,1266) : 0
A
use : 
dir : i
shape : 
(74,866):(294,1124) : 0
VSS
use : g
dir : b
shape : 
(1304,-160):(1400,160) : 0
(1124,-160):(1304,244) : 0
(626,-160):(1124,160) : 0
(446,-160):(626,244) : 0
(0,-160):(446,160) : 0
VDD
use : p
dir : b
shape : 
(1304,2240):(1400,2560) : 0
(1124,2156):(1304,2560) : 0
(634,2240):(1124,2560) : 0
(430,2156):(634,2560) : 0
(0,2240):(430,2560) : 0
CLKBUFX2
--pins(4)
Y
use :  
dir : o
shape : 
(1166,602):(1286,1420) : 0
(1164,550):(1166,1420) : 0
(870,550):(1164,712) : 0
(1124,1254):(1164,1472) : 0
(848,1310):(1124,1472) : 0
A
use : 
dir : i
shape : 
(74,836):(478,1076) : 0
VSS
use : g
dir : b
shape : 
(646,-160):(1400,160) : 0
(466,-160):(646,244) : 0
(0,-160):(466,160) : 0
VDD
use : p
dir : b
shape : 
(626,2240):(1400,2560) : 0
(596,2156):(626,2560) : 0
(474,2130):(596,2560) : 0
(446,2156):(474,2560) : 0
(0,2240):(446,2560) : 0
CLKBUFX20
--pins(4)
Y
use :  
dir : o
shape : 
(7828,572):(7936,1828) : 0
(7114,536):(7828,1828) : 0
(2492,536):(7114,896) : 0
(7074,1266):(7114,1678) : 0
(2472,1318):(7074,1678) : 0
A
use : 
dir : i
shape : 
(1636,948):(1984,1110) : 0
(1514,878):(1636,1110) : 0
(308,948):(1514,1110) : 0
VSS
use : g
dir : b
shape : 
(5728,-160):(8400,160) : 0
(5546,-160):(5728,396) : 0
(5048,-160):(5546,160) : 0
(4868,-160):(5048,396) : 0
(4370,-160):(4868,160) : 0
(4190,-160):(4370,396) : 0
(3690,-160):(4190,160) : 0
(3510,-160):(3690,396) : 0
(3012,-160):(3510,160) : 0
(2832,-160):(3012,396) : 0
(2334,-160):(2832,160) : 0
(2154,-160):(2334,428) : 0
(1570,-160):(2154,160) : 0
(1390,-160):(1570,428) : 0
(806,-160):(1390,160) : 0
(626,-160):(806,428) : 0
(0,-160):(626,160) : 0
VDD
use : p
dir : b
shape : 
(7764,2240):(8400,2560) : 0
(7734,2156):(7764,2560) : 0
(7612,2130):(7734,2560) : 0
(7584,2156):(7612,2560) : 0
(7064,2240):(7584,2560) : 0
(6884,1978):(7064,2560) : 0
(6384,2240):(6884,2560) : 0
(6204,1978):(6384,2560) : 0
(5706,2240):(6204,2560) : 0
(5526,1978):(5706,2560) : 0
(5028,2240):(5526,2560) : 0
(4846,1978):(5028,2560) : 0
(4348,2240):(4846,2560) : 0
(4168,1978):(4348,2560) : 0
(3670,2240):(4168,2560) : 0
(3490,1944):(3670,2560) : 0
(2990,2240):(3490,2560) : 0
(2810,1944):(2990,2560) : 0
(2312,2240):(2810,2560) : 0
(2132,1908):(2312,2560) : 0
(1634,2240):(2132,2560) : 0
(1454,1908):(1634,2560) : 0
(954,2240):(1454,2560) : 0
(774,1908):(954,2560) : 0
(276,2240):(774,2560) : 0
(96,1908):(276,2560) : 0
(0,2240):(96,2560) : 0
CLKBUFX1
--pins(4)
Y
use :  
dir : o
shape : 
(1164,580):(1286,1452) : 0
(1018,580):(1164,690) : 0
(1124,1254):(1164,1452) : 0
(976,1342):(1124,1452) : 0
(838,528):(1018,690) : 0
(796,1342):(976,1504) : 0
A
use : 
dir : i
shape : 
(74,836):(430,1070) : 0
VSS
use : g
dir : b
shape : 
(594,-160):(1400,160) : 0
(414,-160):(594,244) : 0
(0,-160):(414,160) : 0
VDD
use : p
dir : b
shape : 
(626,2240):(1400,2560) : 0
(446,2156):(626,2560) : 0
(0,2240):(446,2560) : 0
CLKBUFX16
--pins(4)
Y
use :  
dir : o
shape : 
(6378,572):(6486,1828) : 0
(5672,536):(6378,1828) : 0
(2136,536):(5672,896) : 0
(5632,1266):(5672,1678) : 0
(2168,1318):(5632,1678) : 0
A
use : 
dir : i
shape : 
(674,852):(1594,1014) : 0
VSS
use : g
dir : b
shape : 
(4778,-160):(6600,160) : 0
(4600,-160):(4778,396) : 0
(4022,-160):(4600,160) : 0
(3842,-160):(4022,396) : 0
(3326,-160):(3842,160) : 0
(3148,-160):(3326,396) : 0
(2652,-160):(3148,160) : 0
(2474,-160):(2652,396) : 0
(1978,-160):(2474,160) : 0
(1800,-160):(1978,396) : 0
(1222,-160):(1800,160) : 0
(1042,-160):(1222,396) : 0
(0,-160):(1042,160) : 0
VDD
use : p
dir : b
shape : 
(6094,2240):(6600,2560) : 0
(5916,1978):(6094,2560) : 0
(5400,2240):(5916,2560) : 0
(5222,1944):(5400,2560) : 0
(4726,2240):(5222,2560) : 0
(4548,1944):(4726,2560) : 0
(4052,2240):(4548,2560) : 0
(3874,1944):(4052,2560) : 0
(3358,2240):(3874,2560) : 0
(3178,1944):(3358,2560) : 0
(2684,2240):(3178,2560) : 0
(2506,1944):(2684,2560) : 0
(2010,2240):(2506,2560) : 0
(1832,1944):(2010,2560) : 0
(1316,2240):(1832,2560) : 0
(1136,1754):(1316,2560) : 0
(622,2240):(1136,2560) : 0
(592,2156):(622,2560) : 0
(472,2130):(592,2560) : 0
(442,2156):(472,2560) : 0
(0,2240):(442,2560) : 0
BUFXL
--pins(4)
Y
use :  
dir : o
shape : 
(1164,548):(1286,1452) : 0
(996,548):(1164,658) : 0
(1124,1254):(1164,1452) : 0
(976,1342):(1124,1452) : 0
(816,496):(996,658) : 0
(796,1342):(976,1504) : 0
A
use : 
dir : i
shape : 
(74,836):(430,1070) : 0
VSS
use : g
dir : b
shape : 
(594,-160):(1400,160) : 0
(414,-160):(594,244) : 0
(0,-160):(414,160) : 0
VDD
use : p
dir : b
shape : 
(626,2240):(1400,2560) : 0
(446,2156):(626,2560) : 0
(0,2240):(446,2560) : 0
BUFX8
--pins(4)
Y
use :  
dir : o
shape : 
(2440,866):(2728,1534) : 0
(2262,866):(2440,1548) : 0
(1894,614):(2262,1548) : 0
(1854,614):(1894,880) : 0
(1854,1252):(1894,1548) : 0
(1218,614):(1854,842) : 0
(1174,1320):(1854,1548) : 0
A
use : 
dir : i
shape : 
(596,948):(744,1110) : 0
(472,878):(596,1110) : 0
(308,948):(472,1110) : 0
VSS
use : g
dir : b
shape : 
(2436,-160):(3200,160) : 0
(2252,-160):(2436,422) : 0
(1746,-160):(2252,160) : 0
(1562,-160):(1746,422) : 0
(1056,-160):(1562,160) : 0
(872,-160):(1056,396) : 0
(280,-160):(872,160) : 0
(96,-160):(280,422) : 0
(0,-160):(96,160) : 0
VDD
use : p
dir : b
shape : 
(2392,2240):(3200,2560) : 0
(2208,1754):(2392,2560) : 0
(1702,2240):(2208,2560) : 0
(1520,1754):(1702,2560) : 0
(1012,2240):(1520,2560) : 0
(830,1794):(1012,2560) : 0
(324,2240):(830,2560) : 0
(140,1794):(324,2560) : 0
(0,2240):(140,2560) : 0
BUFX4
--pins(4)
Y
use :  
dir : o
shape : 
(1200,600):(1364,1466) : 0
(1156,600):(1200,1534) : 0
(1112,600):(1156,824) : 0
(1112,1304):(1156,1534) : 0
(928,438):(1112,824) : 0
(928,1304):(1112,1914) : 0
A
use : 
dir : i
shape : 
(76,866):(436,1140) : 0
VSS
use : g
dir : b
shape : 
(1528,-160):(1800,160) : 0
(1342,-160):(1528,244) : 0
(698,-160):(1342,160) : 0
(512,-160):(698,244) : 0
(0,-160):(512,160) : 0
VDD
use : p
dir : b
shape : 
(1528,2240):(1800,2560) : 0
(1342,1906):(1528,2560) : 0
(698,2240):(1342,2560) : 0
(512,1906):(698,2560) : 0
(0,2240):(512,2560) : 0
BUFX3
--pins(4)
Y
use :  
dir : o
shape : 
(938,574):(996,736) : 0
(938,866):(976,1504) : 0
(816,574):(938,1504) : 0
(796,866):(816,1504) : 0
(774,866):(796,1266) : 0
A
use : 
dir : i
shape : 
(74,866):(294,1124) : 0
VSS
use : g
dir : b
shape : 
(1294,-160):(1400,160) : 0
(1114,-160):(1294,244) : 0
(0,-160):(1114,160) : 0
VDD
use : p
dir : b
shape : 
(572,2240):(1400,2560) : 0
(392,2156):(572,2560) : 0
(0,2240):(392,2560) : 0
BUFX2
--pins(4)
Y
use :  
dir : o
shape : 
(1246,878):(1286,988) : 0
(1124,714):(1246,1420) : 0
(1050,714):(1124,824) : 0
(1028,1310):(1124,1420) : 0
(870,662):(1050,824) : 0
(848,1310):(1028,1472) : 0
A
use : 
dir : i
shape : 
(74,836):(472,1076) : 0
VSS
use : g
dir : b
shape : 
(646,-160):(1400,160) : 0
(466,-160):(646,244) : 0
(0,-160):(466,160) : 0
VDD
use : p
dir : b
shape : 
(626,2240):(1400,2560) : 0
(596,2156):(626,2560) : 0
(474,2130):(596,2560) : 0
(446,2156):(474,2560) : 0
(0,2240):(446,2560) : 0
BUFX20
--pins(4)
Y
use :  
dir : o
shape : 
(4664,536):(5486,1828) : 0
(1814,536):(4664,816) : 0
(4624,1366):(4664,1678) : 0
(1792,1398):(4624,1678) : 0
A
use : 
dir : i
shape : 
(936,948):(1326,1110) : 0
(814,878):(936,1110) : 0
(398,948):(814,1110) : 0
VSS
use : g
dir : b
shape : 
(5070,-160):(5600,160) : 0
(4890,-160):(5070,244) : 0
(4370,-160):(4890,160) : 0
(4190,-160):(4370,396) : 0
(3690,-160):(4190,160) : 0
(3510,-160):(3690,396) : 0
(3012,-160):(3510,160) : 0
(2832,-160):(3012,396) : 0
(2334,-160):(2832,160) : 0
(2154,-160):(2334,396) : 0
(1654,-160):(2154,160) : 0
(1474,-160):(1654,430) : 0
(954,-160):(1474,160) : 0
(774,-160):(954,468) : 0
(276,-160):(774,160) : 0
(96,-160):(276,468) : 0
(0,-160):(96,160) : 0
VDD
use : p
dir : b
shape : 
(5048,2240):(5600,2560) : 0
(5020,2156):(5048,2560) : 0
(4898,2130):(5020,2560) : 0
(4868,2156):(4898,2560) : 0
(4348,2240):(4868,2560) : 0
(4168,1978):(4348,2560) : 0
(3670,2240):(4168,2560) : 0
(3490,1978):(3670,2560) : 0
(2990,2240):(3490,2560) : 0
(2810,1944):(2990,2560) : 0
(2312,2240):(2810,2560) : 0
(2132,1944):(2312,2560) : 0
(1634,2240):(2132,2560) : 0
(1454,1746):(1634,2560) : 0
(954,2240):(1454,2560) : 0
(774,1746):(954,2560) : 0
(276,2240):(774,2560) : 0
(96,1746):(276,2560) : 0
(0,2240):(96,2560) : 0
BUFX1
--pins(4)
Y
use :  
dir : o
shape : 
(1164,548):(1286,1452) : 0
(996,548):(1164,658) : 0
(1124,1254):(1164,1452) : 0
(976,1342):(1124,1452) : 0
(816,496):(996,658) : 0
(796,1342):(976,1504) : 0
A
use : 
dir : i
shape : 
(74,836):(430,1070) : 0
VSS
use : g
dir : b
shape : 
(594,-160):(1400,160) : 0
(414,-160):(594,244) : 0
(0,-160):(414,160) : 0
VDD
use : p
dir : b
shape : 
(626,2240):(1400,2560) : 0
(446,2156):(626,2560) : 0
(0,2240):(446,2560) : 0
BUFX16
--pins(4)
Y
use :  
dir : o
shape : 
(3654,536):(4484,1828) : 0
(1490,536):(3654,816) : 0
(3614,1350):(3654,1678) : 0
(1834,1398):(3614,1678) : 0
A
use : 
dir : i
shape : 
(946,1042):(1094,1204) : 0
(822,1042):(946,1254) : 0
(310,1042):(822,1204) : 0
VSS
use : g
dir : b
shape : 
(4138,-160):(4600,160) : 0
(3956,-160):(4138,244) : 0
(3410,-160):(3956,160) : 0
(3228,-160):(3410,396) : 0
(2702,-160):(3228,160) : 0
(2520,-160):(2702,396) : 0
(2016,-160):(2520,160) : 0
(1834,-160):(2016,396) : 0
(1308,-160):(1834,160) : 0
(1126,-160):(1308,432) : 0
(622,-160):(1126,160) : 0
(440,-160):(622,430) : 0
(0,-160):(440,160) : 0
VDD
use : p
dir : b
shape : 
(4504,2240):(4600,2560) : 0
(4322,2156):(4504,2560) : 0
(3774,2240):(4322,2560) : 0
(3592,2156):(3774,2560) : 0
(3046,2240):(3592,2560) : 0
(2862,1944):(3046,2560) : 0
(2358,2240):(2862,2560) : 0
(2176,1944):(2358,2560) : 0
(1672,2240):(2176,2560) : 0
(1490,1944):(1672,2560) : 0
(966,2240):(1490,2560) : 0
(782,1646):(966,2560) : 0
(278,2240):(782,2560) : 0
(96,1646):(278,2560) : 0
(0,2240):(96,2560) : 0
BUFX12
--pins(4)
Y
use :  
dir : o
shape : 
(2638,600):(3482,1534) : 0
(2596,642):(2638,880) : 0
(2596,1252):(2638,1514) : 0
(1538,642):(2596,804) : 0
(1494,1352):(2596,1514) : 0
A
use : 
dir : i
shape : 
(602,948):(1108,1110) : 0
(478,878):(602,1110) : 0
(388,948):(478,1110) : 0
VSS
use : g
dir : b
shape : 
(3470,-160):(3600,160) : 0
(3284,-160):(3470,422) : 0
(2770,-160):(3284,160) : 0
(2586,-160):(2770,422) : 0
(2072,-160):(2586,160) : 0
(1888,-160):(2072,430) : 0
(1374,-160):(1888,160) : 0
(1190,-160):(1374,430) : 0
(654,-160):(1190,160) : 0
(470,-160):(654,244) : 0
(0,-160):(470,160) : 0
VDD
use : p
dir : b
shape : 
(3502,2240):(3600,2560) : 0
(3316,1944):(3502,2560) : 0
(2754,2240):(3316,2560) : 0
(2570,1944):(2754,2560) : 0
(2030,2240):(2570,2560) : 0
(1844,1944):(2030,2560) : 0
(1330,2240):(1844,2560) : 0
(1146,1794):(1330,2560) : 0
(632,2240):(1146,2560) : 0
(448,1794):(632,2560) : 0
(0,2240):(448,2560) : 0
AOI33X1
--pins(9)
Y
use :  
dir : o
shape : 
(2646,1146):(2686,1254) : 0
(2564,430):(2646,1492) : 0
(2524,430):(2564,1534) : 0
(1072,430):(2524,540) : 0
(2504,1384):(2524,1534) : 0
(2322,1384):(2504,1824) : 0
(1864,1384):(2322,1492) : 0
(1560,1384):(1864,1546) : 0
B2
use : 
dir : i
shape : 
(74,838):(446,1022) : 0
B1
use :  
dir : i
shape : 
(398,1134):(782,1320) : 0
B0
use :  
dir : i
shape : 
(754,790):(1132,1000) : 0
A2
use :  
dir : i
shape : 
(2068,766):(2336,1014) : 0
A1
use :  
dir : i
shape : 
(1866,1134):(2076,1266) : 0
(1686,1092):(1866,1266) : 0
A0
use :  
dir : i
shape : 
(1278,1092):(1552,1266) : 0
(1164,1146):(1278,1254) : 0
VSS
use : g
dir : b
shape : 
(2248,-160):(2800,160) : 0
(2068,-160):(2248,244) : 0
(276,-160):(2068,160) : 0
(96,-160):(276,650) : 0
(0,-160):(96,160) : 0
VDD
use : p
dir : b
shape : 
(1060,2240):(2800,2560) : 0
(880,2156):(1060,2560) : 0
(276,2240):(880,2560) : 0
(96,1464):(276,2560) : 0
(0,2240):(96,2560) : 0
AOI32X4
--pins(8)
Y
use :  
dir : o
shape : 
(3442,866):(3524,1534) : 0
(3316,714):(3442,1534) : 0
(3150,714):(3316,824) : 0
(2954,1304):(3316,1466) : 0
(2964,662):(3150,824) : 0
B1
use : 
dir : i
shape : 
(1956,1134):(2064,1466) : 0
(1828,1036):(1956,1466) : 0
B0
use :  
dir : i
shape : 
(1156,1134):(1434,1408) : 0
A2
use :  
dir : i
shape : 
(76,750):(418,1000) : 0
A1
use :  
dir : i
shape : 
(436,1134):(816,1374) : 0
A0
use :  
dir : i
shape : 
(796,822):(1132,1000) : 0
VSS
use : g
dir : b
shape : 
(3502,-160):(3600,160) : 0
(3316,-160):(3502,424) : 0
(2770,-160):(3316,160) : 0
(2646,-160):(2770,422) : 0
(2008,-160):(2646,160) : 0
(1822,-160):(2008,244) : 0
(284,-160):(1822,160) : 0
(98,-160):(284,550) : 0
(0,-160):(98,160) : 0
VDD
use : p
dir : b
shape : 
(3488,2240):(3600,2560) : 0
(3302,1794):(3488,2560) : 0
(2788,2240):(3302,2560) : 0
(2602,1794):(2788,2560) : 0
(970,2240):(2602,2560) : 0
(786,2156):(970,2560) : 0
(292,2240):(786,2560) : 0
(82,2156):(292,2560) : 0
(0,2240):(82,2560) : 0
AOI32X1
--pins(8)
Y
use :  
dir : o
shape : 
(2350,446):(2480,1640) : 0
(2308,446):(2350,612) : 0
(1722,1530):(2350,1640) : 0
(1136,446):(2308,554) : 0
B1
use : 
dir : i
shape : 
(1754,762):(2108,988) : 0
B0
use :  
dir : i
shape : 
(1424,1120):(1778,1280) : 0
A2
use :  
dir : i
shape : 
(78,800):(450,1000) : 0
A1
use :  
dir : i
shape : 
(492,1142):(832,1360) : 0
A0
use :  
dir : i
shape : 
(822,766):(1194,1000) : 0
VSS
use : g
dir : b
shape : 
(2088,-160):(2600,160) : 0
(1896,-160):(2088,244) : 0
(262,-160):(1896,160) : 0
(132,-160):(262,650) : 0
(0,-160):(132,160) : 0
VDD
use : p
dir : b
shape : 
(1104,2240):(2600,2560) : 0
(912,1850):(1104,2560) : 0
(292,2240):(912,2560) : 0
(102,1600):(292,2560) : 0
(0,2240):(102,2560) : 0
AOI31XL
--pins(7)
Y
use :  
dir : o
shape : 
(1672,560):(1682,722) : 0
(1546,560):(1672,1580) : 0
(1102,560):(1546,670) : 0
B0
use : 
dir : i
shape : 
(1284,1130):(1410,1312) : 0
(1070,1134):(1284,1312) : 0
A2
use :  
dir : i
shape : 
(76,762):(284,1040) : 0
A1
use :  
dir : i
shape : 
(436,1134):(810,1300) : 0
A0
use :  
dir : i
shape : 
(840,780):(1244,1000) : 0
(838,878):(840,988) : 0
VSS
use : g
dir : b
shape : 
(1672,-160):(1800,160) : 0
(1486,-160):(1672,244) : 0
(284,-160):(1486,160) : 0
(98,-160):(284,550) : 0
(0,-160):(98,160) : 0
VDD
use : p
dir : b
shape : 
(1004,2240):(1800,2560) : 0
(818,2156):(1004,2560) : 0
(298,2240):(818,2560) : 0
(96,2156):(298,2560) : 0
(0,2240):(96,2560) : 0
AOI31X1
--pins(7)
Y
use :  
dir : o
shape : 
(1650,402):(1682,1512) : 0
(1558,402):(1650,1916) : 0
(1516,402):(1558,734) : 0
(1524,1402):(1558,1916) : 0
(1102,402):(1516,512) : 0
B0
use : 
dir : i
shape : 
(1430,1002):(1432,1166) : 0
(1216,1002):(1430,1266) : 0
(1156,1134):(1216,1266) : 0
A2
use :  
dir : i
shape : 
(76,840):(284,1142) : 0
A1
use :  
dir : i
shape : 
(436,1116):(706,1336) : 0
A0
use :  
dir : i
shape : 
(796,796):(1058,1000) : 0
VSS
use : g
dir : b
shape : 
(1702,-160):(1800,160) : 0
(1516,-160):(1702,244) : 0
(284,-160):(1516,160) : 0
(98,-160):(284,396) : 0
(0,-160):(98,160) : 0
VDD
use : p
dir : b
shape : 
(982,2240):(1800,2560) : 0
(796,1830):(982,2560) : 0
(284,2240):(796,2560) : 0
(98,1832):(284,2560) : 0
(0,2240):(98,2560) : 0
AOI2BB2X4
--pins(7)
Y
use :  
dir : o
shape : 
(4234,334):(4434,1000) : 0
(1856,538):(4234,648) : 0
(1848,1958):(2490,2066) : 0
(1848,442):(1856,648) : 0
(1728,442):(1848,2066) : 0
(1638,1958):(1728,2066) : 0
B1
use : 
dir : i
shape : 
(4026,1174):(4590,1284) : 0
(3906,876):(4026,1284) : 0
(2660,876):(3906,986) : 0
(2362,876):(2660,988) : 0
(2240,876):(2362,1108) : 0
B0
use :  
dir : i
shape : 
(3128,1134):(3394,1336) : 0
A1N
use :  
dir : i
shape : 
(1126,1412):(1274,1522) : 0
(1006,920):(1126,1984) : 0
(274,1874):(1006,1984) : 0
(250,1788):(274,1984) : 0
(128,1124):(250,1984) : 0
A0N
use :  
dir : i
shape : 
(394,816):(640,1052) : 0
VSS
use : g
dir : b
shape : 
(3726,-160):(5200,160) : 0
(3548,-160):(3726,396) : 0
(2264,-160):(3548,160) : 0
(2086,-160):(2264,396) : 0
(1306,-160):(2086,160) : 0
(1126,-160):(1306,244) : 0
(480,-160):(1126,160) : 0
(302,-160):(480,396) : 0
(0,-160):(302,160) : 0
VDD
use : p
dir : b
shape : 
(4506,2240):(5200,2560) : 0
(4328,1960):(4506,2560) : 0
(3834,2240):(4328,2560) : 0
(3656,1960):(3834,2560) : 0
(3162,2240):(3656,2560) : 0
(2984,1960):(3162,2560) : 0
(1450,2240):(2984,2560) : 0
(1272,2156):(1450,2560) : 0
(274,2240):(1272,2560) : 0
(94,2156):(274,2560) : 0
(0,2240):(94,2560) : 0
AOI2BB2X2
--pins(7)
Y
use :  
dir : o
shape : 
(3016,612):(3084,722) : 0
(2892,384):(3016,1954) : 0
(1546,384):(2892,492) : 0
(2608,1846):(2892,1954) : 0
(2406,1846):(2608,2080) : 0
(2374,1934):(2406,2080) : 0
(2188,1972):(2374,2080) : 0
B1
use : 
dir : i
shape : 
(2208,1086):(2402,1474) : 0
(1024,1364):(2208,1474) : 0
B0
use :  
dir : i
shape : 
(2588,758):(2742,996) : 0
(1344,758):(2588,866) : 0
A1N
use :  
dir : i
shape : 
(686,776):(992,1000) : 0
A0N
use :  
dir : i
shape : 
(76,890):(280,1266) : 0
VSS
use : g
dir : b
shape : 
(2144,-160):(3200,160) : 0
(1960,-160):(2144,244) : 0
(1032,-160):(1960,160) : 0
(848,-160):(1032,578) : 0
(280,-160):(848,160) : 0
(96,-160):(280,244) : 0
(0,-160):(96,160) : 0
VDD
use : p
dir : b
shape : 
(3082,2240):(3200,2560) : 0
(2898,2156):(3082,2560) : 0
(1680,2240):(2898,2560) : 0
(1498,1976):(1680,2560) : 0
(992,2240):(1498,2560) : 0
(808,1976):(992,2560) : 0
(0,2240):(808,2560) : 0
AOI2BB2X1
--pins(7)
Y
use :  
dir : o
shape : 
(2194,530):(2324,2098) : 0
(1520,530):(2194,640) : 0
(1978,1134):(2194,1266) : 0
B1
use : 
dir : i
shape : 
(1100,1322):(1406,1534) : 0
B0
use :  
dir : i
shape : 
(1606,1072):(1736,1254) : 0
(1474,1072):(1606,1180) : 0
(1346,1002):(1474,1180) : 0
A1N
use :  
dir : i
shape : 
(106,866):(268,1240) : 0
A0N
use :  
dir : i
shape : 
(448,1072):(696,1302) : 0
VSS
use : g
dir : b
shape : 
(2138,-160):(2600,160) : 0
(1948,-160):(2138,244) : 0
(968,-160):(1948,160) : 0
(776,-160):(968,244) : 0
(292,-160):(776,160) : 0
(102,-160):(292,244) : 0
(0,-160):(102,160) : 0
VDD
use : p
dir : b
shape : 
(1632,2240):(2600,2560) : 0
(1440,1978):(1632,2560) : 0
(292,2240):(1440,2560) : 0
(102,2156):(292,2560) : 0
(0,2240):(102,2560) : 0
AOI2BB1XL
--pins(6)
Y
use :  
dir : o
shape : 
(1584,1678):(1682,1788) : 0
(1460,772):(1584,1814) : 0
(1148,772):(1460,880) : 0
(1022,696):(1148,880) : 0
B0
use : 
dir : i
shape : 
(796,1272):(1064,1534) : 0
A1N
use :  
dir : i
shape : 
(294,1076):(602,1254) : 0
A0N
use :  
dir : i
shape : 
(96,1378):(398,1578) : 0
VSS
use : g
dir : b
shape : 
(692,-160):(1800,160) : 0
(508,-160):(692,244) : 0
(0,-160):(508,160) : 0
VDD
use : p
dir : b
shape : 
(894,2240):(1800,2560) : 0
(710,2156):(894,2560) : 0
(0,2240):(710,2560) : 0
AOI2BB1X1
--pins(6)
Y
use :  
dir : o
shape : 
(1588,584):(1682,1522) : 0
(1558,584):(1588,1972) : 0
(1140,584):(1558,692) : 0
(1462,1412):(1558,1972) : 0
B0
use : 
dir : i
shape : 
(1070,1330):(1072,1522) : 0
(718,1330):(1070,1534) : 0
A1N
use :  
dir : i
shape : 
(300,848):(644,1010) : 0
A0N
use :  
dir : i
shape : 
(76,1134):(436,1358) : 0
VSS
use : g
dir : b
shape : 
(692,-160):(1800,160) : 0
(508,-160):(692,244) : 0
(0,-160):(508,160) : 0
VDD
use : p
dir : b
shape : 
(894,2240):(1800,2560) : 0
(710,2156):(894,2560) : 0
(0,2240):(710,2560) : 0
AOI22XL
--pins(7)
Y
use :  
dir : o
shape : 
(1598,564):(1724,1630) : 0
(1558,564):(1598,722) : 0
(1330,1522):(1598,1630) : 0
(1004,564):(1558,674) : 0
(1146,1496):(1330,1658) : 0
(818,538):(1004,700) : 0
B1
use : 
dir : i
shape : 
(76,792):(338,1022) : 0
B0
use :  
dir : i
shape : 
(650,1120):(834,1298) : 0
(436,1134):(650,1298) : 0
A1
use :  
dir : i
shape : 
(1432,1142):(1462,1304) : 0
(1134,1124):(1432,1304) : 0
A0
use :  
dir : i
shape : 
(1202,850):(1206,1000) : 0
(962,824):(1202,1000) : 0
(834,850):(962,1000) : 0
VSS
use : g
dir : b
shape : 
(1680,-160):(1800,160) : 0
(1494,-160):(1680,244) : 0
(284,-160):(1494,160) : 0
(98,-160):(284,244) : 0
(0,-160):(98,160) : 0
VDD
use : p
dir : b
shape : 
(352,2240):(1800,2560) : 0
(126,2156):(352,2560) : 0
(0,2240):(126,2560) : 0
AOI22X4
--pins(7)
Y
use :  
dir : o
shape : 
(4568,878):(4692,1970) : 0
(4526,600):(4568,1266) : 0
(4048,1860):(4568,1970) : 0
(4362,574):(4526,1266) : 0
(98,574):(4362,684) : 0
(3878,1860):(4048,2066) : 0
(3810,1934):(3878,2066) : 0
(2522,1958):(3810,2066) : 0
B1
use : 
dir : i
shape : 
(2132,876):(2162,986) : 0
(2008,876):(2132,988) : 0
(474,878):(2008,988) : 0
B0
use :  
dir : i
shape : 
(1312,1174):(1540,1284) : 0
(1188,1146):(1312,1284) : 0
(228,1174):(1188,1284) : 0
A1
use :  
dir : i
shape : 
(2576,878):(3744,988) : 0
(2494,878):(2576,1000) : 0
(2370,878):(2494,1308) : 0
A0
use :  
dir : i
shape : 
(4086,1008):(4210,1254) : 0
(2740,1146):(4086,1254) : 0
VSS
use : g
dir : b
shape : 
(3744,-160):(5000,160) : 0
(3560,-160):(3744,406) : 0
(2360,-160):(3560,160) : 0
(2176,-160):(2360,406) : 0
(974,-160):(2176,160) : 0
(790,-160):(974,406) : 0
(0,-160):(790,160) : 0
VDD
use : p
dir : b
shape : 
(2012,2240):(5000,2560) : 0
(1830,1960):(2012,2560) : 0
(1320,2240):(1830,2560) : 0
(1136,1960):(1320,2560) : 0
(628,2240):(1136,2560) : 0
(444,1960):(628,2560) : 0
(0,2240):(444,2560) : 0
AOI22X2
--pins(7)
Y
use :  
dir : o
shape : 
(2960,642):(3084,1522) : 0
(786,642):(2960,752) : 0
(2736,1412):(2960,1522) : 0
(2604,1412):(2736,1578) : 0
(1864,1470):(2604,1578) : 0
B1
use : 
dir : i
shape : 
(1306,912):(1430,1150) : 0
(596,912):(1306,1022) : 0
(492,878):(596,1022) : 0
(370,878):(492,1124) : 0
(226,986):(370,1124) : 0
B0
use :  
dir : i
shape : 
(658,1146):(950,1326) : 0
A1
use :  
dir : i
shape : 
(2712,876):(2836,1102) : 0
(2018,876):(2712,986) : 0
(1888,876):(2018,988) : 0
(1764,876):(1888,1328) : 0
A0
use :  
dir : i
shape : 
(2122,1134):(2414,1322) : 0
VSS
use : g
dir : b
shape : 
(2888,-160):(3200,160) : 0
(2704,-160):(2888,244) : 0
(1574,-160):(2704,160) : 0
(1390,-160):(1574,244) : 0
(280,-160):(1390,160) : 0
(96,-160):(280,610) : 0
(0,-160):(96,160) : 0
VDD
use : p
dir : b
shape : 
(1314,2240):(3200,2560) : 0
(1132,1776):(1314,2560) : 0
(624,2240):(1132,2560) : 0
(442,1776):(624,2560) : 0
(0,2240):(442,2560) : 0
AOI22X1
--pins(7)
Y
use :  
dir : o
shape : 
(1598,530):(1724,1508) : 0
(1558,530):(1598,722) : 0
(1352,1398):(1598,1508) : 0
(982,530):(1558,640) : 0
(1168,1398):(1352,1560) : 0
(796,504):(982,666) : 0
B1
use : 
dir : i
shape : 
(104,842):(290,1178) : 0
B0
use :  
dir : i
shape : 
(478,1134):(830,1326) : 0
A1
use :  
dir : i
shape : 
(1154,1076):(1462,1266) : 0
A0
use :  
dir : i
shape : 
(998,788):(1184,950) : 0
(962,814):(998,950) : 0
(838,814):(962,988) : 0
VSS
use : g
dir : b
shape : 
(1702,-160):(1800,160) : 0
(1516,-160):(1702,244) : 0
(284,-160):(1516,160) : 0
(98,-160):(284,660) : 0
(0,-160):(98,160) : 0
VDD
use : p
dir : b
shape : 
(644,2240):(1800,2560) : 0
(458,2156):(644,2560) : 0
(0,2240):(458,2560) : 0
AOI222XL
--pins(9)
Y
use :  
dir : o
shape : 
(2564,540):(2686,1474) : 0
(96,540):(2564,650) : 0
(2524,1254):(2564,1474) : 0
(2102,1364):(2524,1474) : 0
C1
use :  
dir : i
shape : 
(424,1136):(674,1374) : 0
C0
use :  
dir : i
shape : 
(74,866):(276,1128) : 0
B1
use :  
dir : i
shape : 
(808,822):(1100,1000) : 0
B0
use :  
dir : i
shape : 
(1376,866):(1668,1048) : 0
A1
use :  
dir : i
shape : 
(2212,878):(2396,1210) : 0
A0
use :  
dir : i
shape : 
(1842,784):(2044,1046) : 0
VSS
use : g
dir : b
shape : 
(2572,-160):(2800,160) : 0
(2392,-160):(2572,244) : 0
(1000,-160):(2392,160) : 0
(820,-160):(1000,400) : 0
(0,-160):(820,160) : 0
VDD
use : p
dir : b
shape : 
(616,2240):(2800,2560) : 0
(434,2130):(616,2560) : 0
(0,2240):(434,2560) : 0
AOI222X1
--pins(9)
Y
use :  
dir : o
shape : 
(2564,562):(2686,1486) : 0
(96,562):(2564,672) : 0
(2166,1376):(2564,1486) : 0
C1
use :  
dir : i
shape : 
(464,810):(760,1014) : 0
C0
use :  
dir : i
shape : 
(74,878):(244,1266) : 0
B1
use :  
dir : i
shape : 
(976,1012):(1172,1254) : 0
(814,1146):(976,1254) : 0
B0
use :  
dir : i
shape : 
(1402,866):(1676,1070) : 0
A1
use :  
dir : i
shape : 
(2174,866):(2376,1174) : 0
A0
use :  
dir : i
shape : 
(1824,888):(2026,1254) : 0
VSS
use : g
dir : b
shape : 
(2538,-160):(2800,160) : 0
(2358,-160):(2538,244) : 0
(1016,-160):(2358,160) : 0
(836,-160):(1016,244) : 0
(0,-160):(836,160) : 0
VDD
use : p
dir : b
shape : 
(954,2240):(2800,2560) : 0
(774,1834):(954,2560) : 0
(276,2240):(774,2560) : 0
(96,1882):(276,2560) : 0
(0,2240):(96,2560) : 0
AOI221XL
--pins(8)
Y
use :  
dir : o
shape : 
(2350,472):(2480,1486) : 0
(2308,472):(2350,612) : 0
(2184,1376):(2350,1486) : 0
(1224,472):(2308,580) : 0
(1094,322):(1224,580) : 0
(994,322):(1094,466) : 0
(822,322):(994,430) : 0
C0
use :  
dir : i
shape : 
(2038,1146):(2108,1254) : 0
(1908,866):(2038,1254) : 0
B1
use :  
dir : i
shape : 
(78,626):(292,1000) : 0
B0
use :  
dir : i
shape : 
(450,1124):(754,1342) : 0
A1
use :  
dir : i
shape : 
(1444,748):(1736,988) : 0
A0
use :  
dir : i
shape : 
(976,878):(1106,1226) : 0
(864,878):(976,988) : 0
VSS
use : g
dir : b
shape : 
(1756,-160):(2600,160) : 0
(1564,-160):(1756,244) : 0
(292,-160):(1564,160) : 0
(102,-160):(292,396) : 0
(0,-160):(102,160) : 0
VDD
use : p
dir : b
shape : 
(922,2240):(2600,2560) : 0
(732,2156):(922,2560) : 0
(292,2240):(732,2560) : 0
(102,2156):(292,2560) : 0
(0,2240):(102,2560) : 0
AOI221X2
--pins(8)
Y
use :  
dir : o
shape : 
(3614,624):(3736,1672) : 0
(2914,624):(3614,734) : 0
(3522,1510):(3614,1672) : 0
(2782,600):(2914,734) : 0
(2660,450):(2782,734) : 0
(774,450):(2660,560) : 0
C0
use :  
dir : i
shape : 
(3356,878):(3478,1086) : 0
(2914,878):(3356,988) : 0
B1
use :  
dir : i
shape : 
(1326,986):(1422,1116) : 0
(1124,866):(1326,1116) : 0
(154,1008):(1124,1116) : 0
B0
use :  
dir : i
shape : 
(626,750):(828,860) : 0
(424,612):(626,860) : 0
A1
use :  
dir : i
shape : 
(1986,1190):(3144,1300) : 0
(1864,1146):(1986,1300) : 0
(1834,1190):(1864,1300) : 0
A0
use :  
dir : i
shape : 
(2174,792):(2466,1000) : 0
VSS
use : g
dir : b
shape : 
(3272,-160):(4200,160) : 0
(3092,-160):(3272,396) : 0
(1740,-160):(3092,160) : 0
(1560,-160):(1740,244) : 0
(276,-160):(1560,160) : 0
(96,-160):(276,396) : 0
(0,-160):(96,160) : 0
VDD
use : p
dir : b
shape : 
(1634,2240):(4200,2560) : 0
(1454,1806):(1634,2560) : 0
(954,2240):(1454,2560) : 0
(774,1806):(954,2560) : 0
(276,2240):(774,2560) : 0
(96,1806):(276,2560) : 0
(0,2240):(96,2560) : 0
AOI221X1
--pins(8)
Y
use :  
dir : o
shape : 
(2350,514):(2480,1522) : 0
(1406,514):(2350,624) : 0
(2330,1254):(2350,1508) : 0
(1392,454):(1406,624) : 0
(1264,378):(1392,624) : 0
(822,378):(1264,488) : 0
C0
use :  
dir : i
shape : 
(2088,1146):(2108,1254) : 0
(1958,786):(2088,1254) : 0
B1
use :  
dir : i
shape : 
(98,612):(292,922) : 0
B0
use :  
dir : i
shape : 
(450,1040):(760,1266) : 0
A1
use :  
dir : i
shape : 
(1606,758):(1736,988) : 0
(1334,758):(1606,866) : 0
A0
use :  
dir : i
shape : 
(864,612):(1120,862) : 0
VSS
use : g
dir : b
shape : 
(1756,-160):(2600,160) : 0
(1564,-160):(1756,244) : 0
(292,-160):(1564,160) : 0
(102,-160):(292,458) : 0
(0,-160):(102,160) : 0
VDD
use : p
dir : b
shape : 
(1012,2240):(2600,2560) : 0
(822,1832):(1012,2560) : 0
(292,2240):(822,2560) : 0
(102,1832):(292,2560) : 0
(0,2240):(102,2560) : 0
AOI21XL
--pins(6)
Y
use :  
dir : o
shape : 
(1268,590):(1286,1254) : 0
(1164,590):(1268,1660) : 0
(774,590):(1164,700) : 0
(1146,1146):(1164,1660) : 0
B0
use :  
dir : i
shape : 
(724,822):(1026,1000) : 0
A1
use :  
dir : i
shape : 
(90,834):(276,1124) : 0
A0
use :  
dir : i
shape : 
(424,1134):(758,1324) : 0
VSS
use : g
dir : b
shape : 
(1252,-160):(1400,160) : 0
(1072,-160):(1252,244) : 0
(276,-160):(1072,160) : 0
(96,-160):(276,662) : 0
(0,-160):(96,160) : 0
VDD
use : p
dir : b
shape : 
(626,2240):(1400,2560) : 0
(446,2156):(626,2560) : 0
(0,2240):(446,2560) : 0
AOI21X4
--pins(6)
Y
use :  
dir : o
shape : 
(3336,1792):(3426,1954) : 0
(3240,1158):(3336,1954) : 0
(3210,1158):(3240,1928) : 0
(3164,1158):(3210,1266) : 0
(2728,1820):(3210,1928) : 0
(2956,600):(3164,1266) : 0
(2638,674):(2956,784) : 0
(2542,1792):(2728,1954) : 0
(2416,548):(2638,784) : 0
(98,548):(2416,658) : 0
B0
use :  
dir : i
shape : 
(2476,992):(2804,1270) : 0
A1
use :  
dir : i
shape : 
(2136,904):(2196,1066) : 0
(2010,784):(2136,1066) : 0
(1322,784):(2010,892) : 0
(984,784):(1322,988) : 0
(830,784):(984,1014) : 0
(800,852):(830,1014) : 0
A0
use :  
dir : i
shape : 
(1614,1146):(1682,1254) : 0
(1490,1060):(1614,1254) : 0
(436,1140):(1490,1250) : 0
(414,1134):(436,1250) : 0
(290,938):(414,1250) : 0
(230,938):(290,1148) : 0
VSS
use : g
dir : b
shape : 
(3100,-160):(3600,160) : 0
(2916,-160):(3100,244) : 0
(2380,-160):(2916,160) : 0
(2196,-160):(2380,396) : 0
(984,-160):(2196,160) : 0
(800,-160):(984,396) : 0
(0,-160):(800,160) : 0
VDD
use : p
dir : b
shape : 
(2030,2240):(3600,2560) : 0
(1844,1882):(2030,2560) : 0
(1330,2240):(1844,2560) : 0
(1146,1882):(1330,2560) : 0
(632,2240):(1146,2560) : 0
(448,1882):(632,2560) : 0
(0,2240):(448,2560) : 0
AOI21X2
--pins(6)
Y
use :  
dir : o
shape : 
(2060,690):(2190,1578) : 0
(1734,690):(2060,800) : 0
(1978,1412):(2060,1578) : 0
(1948,1470):(1978,1578) : 0
(1542,536):(1734,800) : 0
(600,690):(1542,800) : 0
(470,588):(600,800) : 0
(292,588):(470,698) : 0
(102,536):(292,698) : 0
B0
use :  
dir : i
shape : 
(1660,970):(1872,1254) : 0
(1606,1146):(1660,1254) : 0
A1
use :  
dir : i
shape : 
(622,1190):(1036,1338) : 0
(492,1146):(622,1338) : 0
A0
use :  
dir : i
shape : 
(292,914):(1526,1024) : 0
(78,866):(292,1060) : 0
VSS
use : g
dir : b
shape : 
(2164,-160):(2600,160) : 0
(1972,-160):(2164,244) : 0
(1012,-160):(1972,160) : 0
(822,-160):(1012,550) : 0
(0,-160):(822,160) : 0
VDD
use : p
dir : b
shape : 
(1374,2240):(2600,2560) : 0
(1182,1776):(1374,2560) : 0
(652,2240):(1182,2560) : 0
(462,1776):(652,2560) : 0
(0,2240):(462,2560) : 0
AOI21X1
--pins(6)
Y
use :  
dir : o
shape : 
(1206,642):(1328,1880) : 0
(954,642):(1206,752) : 0
(1164,1412):(1206,1880) : 0
(1114,1720):(1164,1880) : 0
(774,590):(954,752) : 0
B0
use :  
dir : i
shape : 
(954,878):(1084,1254) : 0
(814,878):(954,988) : 0
A1
use :  
dir : i
shape : 
(276,984):(282,1230) : 0
(100,866):(276,1230) : 0
A0
use :  
dir : i
shape : 
(586,1136):(758,1246) : 0
(464,612):(586,1246) : 0
VSS
use : g
dir : b
shape : 
(1252,-160):(1400,160) : 0
(1072,-160):(1252,244) : 0
(276,-160):(1072,160) : 0
(96,-160):(276,668) : 0
(0,-160):(96,160) : 0
VDD
use : p
dir : b
shape : 
(616,2240):(1400,2560) : 0
(434,1704):(616,2560) : 0
(0,2240):(434,2560) : 0
AND4X4
--pins(7)
Y
use :  
dir : o
shape : 
(3518,1134):(3560,1800) : 0
(3392,712):(3518,1800) : 0
(3352,662):(3392,1800) : 0
(3350,662):(3352,878) : 0
(3350,1134):(3352,1800) : 0
(3140,662):(3350,824) : 0
(3064,1630):(3350,1800) : 0
(2876,1630):(3064,2078) : 0
D
use :  
dir : i
shape : 
(2656,878):(2728,988) : 0
(2528,878):(2656,1300) : 0
(2426,1134):(2528,1300) : 0
(2356,1190):(2426,1300) : 0
(2228,1190):(2356,1776) : 0
(290,1666):(2228,1776) : 0
(290,1280):(292,1534) : 0
(162,1280):(290,1776) : 0
(78,1280):(162,1534) : 0
C
use :  
dir : i
shape : 
(1976,758):(2102,1442) : 0
(1896,758):(1976,878) : 0
(688,758):(1896,866) : 0
(688,1078):(728,1272) : 0
(562,758):(688,1272) : 0
(440,986):(562,1272) : 0
B
use :  
dir : i
shape : 
(1532,978):(1742,1258) : 0
(920,978):(1532,1088) : 0
A
use :  
dir : i
shape : 
(1158,1250):(1378,1546) : 0
VSS
use : g
dir : b
shape : 
(3724,-160):(4000,160) : 0
(3538,-160):(3724,422) : 0
(2932,-160):(3538,160) : 0
(2744,-160):(2932,500) : 0
(286,-160):(2744,160) : 0
(100,-160):(286,668) : 0
(0,-160):(100,160) : 0
VDD
use : p
dir : b
shape : 
(3502,2240):(4000,2560) : 0
(3286,2156):(3502,2560) : 0
(2450,2240):(3286,2560) : 0
(2262,2156):(2450,2560) : 0
(1564,2240):(2262,2560) : 0
(1378,2156):(1564,2560) : 0
(716,2240):(1378,2560) : 0
(502,2156):(716,2560) : 0
(0,2240):(502,2560) : 0
AND4X2
--pins(7)
Y
use :  
dir : o
shape : 
(2098,1400):(2122,1534) : 0
(2062,716):(2098,1534) : 0
(1970,398):(2062,1928) : 0
(1934,398):(1970,826) : 0
(1934,1296):(1970,1928) : 0
D
use :  
dir : i
shape : 
(1388,1048):(1466,1212) : 0
(1220,878):(1388,1212) : 0
C
use :  
dir : i
shape : 
(956,1162):(1084,1522) : 0
(852,1412):(956,1522) : 0
B
use :  
dir : i
shape : 
(558,1074):(716,1292) : 0
(444,1074):(558,1290) : 0
A
use :  
dir : i
shape : 
(78,796):(314,1112) : 0
VSS
use : g
dir : b
shape : 
(1630,-160):(2200,160) : 0
(1442,-160):(1630,244) : 0
(0,-160):(1442,160) : 0
VDD
use : p
dir : b
shape : 
(1676,2240):(2200,2560) : 0
(1448,2128):(1676,2560) : 0
(1028,2240):(1448,2560) : 0
(838,2156):(1028,2560) : 0
(316,2240):(838,2560) : 0
(98,2156):(316,2560) : 0
(0,2240):(98,2560) : 0
AND4X1
--pins(7)
Y
use :  
dir : o
shape : 
(2088,1522):(2122,1810) : 0
(1962,488):(2088,1810) : 0
(1900,488):(1962,650) : 0
(1912,1522):(1962,1810) : 0
(1900,1600):(1912,1810) : 0
D
use :  
dir : i
shape : 
(1406,1146):(1714,1392) : 0
C
use :  
dir : i
shape : 
(784,1134):(1022,1392) : 0
B
use :  
dir : i
shape : 
(350,798):(656,1090) : 0
A
use :  
dir : i
shape : 
(78,1230):(294,1552) : 0
VSS
use : g
dir : b
shape : 
(1666,-160):(2200,160) : 0
(1478,-160):(1666,244) : 0
(0,-160):(1478,160) : 0
VDD
use : p
dir : b
shape : 
(1722,2240):(2200,2560) : 0
(516,2156):(1722,2560) : 0
(0,2240):(516,2560) : 0
AOI211XL
--pins(7)
Y
use :  
dir : o
shape : 
(1598,548):(1724,1522) : 0
(796,548):(1598,658) : 0
(1516,1412):(1598,1522) : 0
C0
use :  
dir : i
shape : 
(824,1110):(1160,1290) : 0
B0
use :  
dir : i
shape : 
(1348,866):(1472,1184) : 0
(1154,866):(1348,1000) : 0
A1
use :  
dir : i
shape : 
(76,930):(284,1266) : 0
A0
use :  
dir : i
shape : 
(434,786):(750,1000) : 0
VSS
use : g
dir : b
shape : 
(1342,-160):(1800,160) : 0
(1156,-160):(1342,244) : 0
(284,-160):(1156,160) : 0
(98,-160):(284,560) : 0
(0,-160):(98,160) : 0
VDD
use : p
dir : b
shape : 
(590,2240):(1800,2560) : 0
(404,2156):(590,2560) : 0
(0,2240):(404,2560) : 0
AOI211X2
--pins(7)
Y
use :  
dir : o
shape : 
(2942,498):(3066,1522) : 0
(2828,498):(2942,608) : 0
(2354,1412):(2942,1522) : 0
(2646,446):(2828,608) : 0
(1960,472):(2646,580) : 0
(2200,1412):(2354,1614) : 0
(2172,1452):(2200,1614) : 0
(1524,446):(1960,608) : 0
(1498,446):(1524,580) : 0
(286,472):(1498,580) : 0
(102,446):(286,608) : 0
C0
use :  
dir : i
shape : 
(2690,730):(2814,1078) : 0
(2564,730):(2690,878) : 0
(1810,730):(2564,840) : 0
(1686,730):(1810,1254) : 0
(1538,1100):(1686,1254) : 0
B0
use :  
dir : i
shape : 
(2042,1100):(2414,1290) : 0
A1
use :  
dir : i
shape : 
(472,1078):(798,1254) : 0
A0
use :  
dir : i
shape : 
(1202,988):(1230,1242) : 0
(1078,798):(1202,1242) : 0
(414,798):(1078,908) : 0
(1048,1080):(1078,1242) : 0
(240,772):(414,934) : 0
(232,772):(240,988) : 0
(116,798):(232,988) : 0
VSS
use : g
dir : b
shape : 
(2416,-160):(3200,160) : 0
(2232,-160):(2416,244) : 0
(996,-160):(2232,160) : 0
(814,-160):(996,244) : 0
(0,-160):(814,160) : 0
VDD
use : p
dir : b
shape : 
(1318,2240):(3200,2560) : 0
(1134,1850):(1318,2560) : 0
(628,2240):(1134,2560) : 0
(444,1850):(628,2560) : 0
(0,2240):(444,2560) : 0
AOI211X1
--pins(7)
Y
use :  
dir : o
shape : 
(1680,522):(1734,1522) : 0
(1642,522):(1680,1950) : 0
(1610,384):(1642,1950) : 0
(1516,384):(1610,684) : 0
(1494,1322):(1610,1950) : 0
(1000,384):(1516,492) : 0
(876,384):(1000,658) : 0
(796,548):(876,658) : 0
C0
use :  
dir : i
shape : 
(796,1030):(1116,1266) : 0
B0
use :  
dir : i
shape : 
(1370,872):(1484,1072) : 0
(1358,872):(1370,1522) : 0
(1244,962):(1358,1522) : 0
(1198,1412):(1244,1522) : 0
A1
use :  
dir : i
shape : 
(76,1048):(352,1290) : 0
A0
use :  
dir : i
shape : 
(644,800):(780,910) : 0
(478,612):(644,910) : 0
VSS
use : g
dir : b
shape : 
(1280,-160):(1800,160) : 0
(1094,-160):(1280,244) : 0
(284,-160):(1094,160) : 0
(98,-160):(284,520) : 0
(0,-160):(98,160) : 0
VDD
use : p
dir : b
shape : 
(632,2240):(1800,2560) : 0
(448,1818):(632,2560) : 0
(0,2240):(448,2560) : 0
AND3X1
--pins(6)
Y
use :  
dir : o
shape : 
(1592,548):(1718,1978) : 0
(1468,548):(1592,710) : 0
(1516,1658):(1592,1978) : 0
C
use :  
dir : i
shape : 
(794,816):(1078,1022) : 0
B
use :  
dir : i
shape : 
(368,1354):(644,1572) : 0
A
use :  
dir : i
shape : 
(76,852):(316,1096) : 0
VSS
use : g
dir : b
shape : 
(1276,-160):(1800,160) : 0
(1090,-160):(1276,244) : 0
(0,-160):(1090,160) : 0
VDD
use : p
dir : b
shape : 
(1388,2240):(1800,2560) : 0
(1388,1342):(1468,1444) : 0
(1262,1342):(1388,2560) : 0
(720,2240):(1262,2560) : 0
(718,2156):(720,2560) : 0
(540,2130):(718,2560) : 0
(534,2156):(540,2560) : 0
(0,2240):(534,2560) : 0
AND2XL
--pins(5)
Y
use :  
dir : o
shape : 
(1248,1134):(1326,1266) : 0
(1126,688):(1248,1690) : 0
B
use :  
dir : i
shape : 
(438,1128):(640,1404) : 0
A
use :  
dir : i
shape : 
(80,866):(300,1102) : 0
VSS
use : g
dir : b
shape : 
(950,-160):(1400,160) : 0
(768,-160):(950,244) : 0
(0,-160):(768,160) : 0
VDD
use : p
dir : b
shape : 
(742,2240):(1400,2560) : 0
(244,2156):(742,2560) : 0
(0,2240):(244,2560) : 0
AND2X4
--pins(5)
Y
use :  
dir : o
shape : 
(1720,866):(1724,1534) : 0
(1568,662):(1720,1596) : 0
(1516,652):(1568,1596) : 0
(1184,652):(1516,866) : 0
(1160,1434):(1516,1596) : 0
B
use :  
dir : i
shape : 
(644,942):(750,1124) : 0
(624,942):(644,1572) : 0
(518,1014):(624,1572) : 0
(436,1254):(518,1572) : 0
A
use :  
dir : i
shape : 
(284,964):(290,1148) : 0
(76,964):(284,1320) : 0
VSS
use : g
dir : b
shape : 
(1696,-160):(1800,160) : 0
(1510,-160):(1696,486) : 0
(960,-160):(1510,160) : 0
(774,-160):(960,244) : 0
(0,-160):(774,160) : 0
VDD
use : p
dir : b
shape : 
(1696,2240):(1800,2560) : 0
(1510,1828):(1696,2560) : 0
(974,2240):(1510,2560) : 0
(788,2156):(974,2560) : 0
(292,2240):(788,2560) : 0
(92,2156):(292,2560) : 0
(0,2240):(92,2560) : 0
AND2X2
--pins(5)
Y
use :  
dir : o
shape : 
(1284,454):(1308,1534) : 0
(1186,390):(1284,2004) : 0
(1164,390):(1186,878) : 0
(1104,1376):(1186,2004) : 0
(1104,390):(1164,780) : 0
B
use :  
dir : i
shape : 
(424,1666):(722,1870) : 0
A
use :  
dir : i
shape : 
(276,1008):(404,1170) : 0
(74,1008):(276,1266) : 0
VSS
use : g
dir : b
shape : 
(880,-160):(1400,160) : 0
(700,-160):(880,244) : 0
(0,-160):(700,160) : 0
VDD
use : p
dir : b
shape : 
(302,2240):(1400,2560) : 0
(96,2156):(302,2560) : 0
(0,2240):(96,2560) : 0
AND2X1
--pins(5)
Y
use :  
dir : o
shape : 
(1248,1134):(1326,1266) : 0
(1248,640):(1278,878) : 0
(1248,1464):(1278,1854) : 0
(1126,640):(1248,1854) : 0
(1124,640):(1126,878) : 0
(1098,1464):(1126,1854) : 0
(1098,640):(1124,802) : 0
B
use :  
dir : i
shape : 
(424,1102):(644,1378) : 0
A
use :  
dir : i
shape : 
(80,866):(300,1102) : 0
VSS
use : g
dir : b
shape : 
(950,-160):(1400,160) : 0
(768,-160):(950,244) : 0
(0,-160):(768,160) : 0
VDD
use : p
dir : b
shape : 
(930,2240):(1400,2560) : 0
(694,2156):(930,2560) : 0
(418,2240):(694,2560) : 0
(238,2156):(418,2560) : 0
(0,2240):(238,2560) : 0
ADDHXL
--pins(6)
S
use :  
dir : o
shape : 
(2400,1412):(2426,1526) : 0
(2272,774):(2400,1526) : 0
(1922,774):(2272,884) : 0
(1878,1416):(2272,1526) : 0
(1796,522):(1922,884) : 0
(1752,1416):(1878,1754) : 0
CO
use :  
dir : o
shape : 
(3870,878):(3882,988) : 0
(3744,300):(3870,1830) : 0
(3582,1722):(3744,1830) : 0
B
use :  
dir : i
shape : 
(1626,1872):(3166,1980) : 0
(1986,1016):(2112,1304) : 0
(1626,1196):(1986,1304) : 0
(1498,1196):(1626,1980) : 0
(1168,1364):(1498,1534) : 0
(978,1364):(1168,1474) : 0
A
use :  
dir : i
shape : 
(2854,1100):(3196,1300) : 0
VSS
use : g
dir : b
shape : 
(3504,-160):(4000,160) : 0
(3316,-160):(3504,432) : 0
(2790,-160):(3316,160) : 0
(2604,-160):(2790,244) : 0
(706,-160):(2604,160) : 0
(518,-160):(706,244) : 0
(0,-160):(518,160) : 0
VDD
use : p
dir : b
shape : 
(3458,2240):(4000,2560) : 0
(3270,2156):(3458,2560) : 0
(2614,2240):(3270,2560) : 0
(2426,2156):(2614,2560) : 0
(706,2240):(2426,2560) : 0
(518,2156):(706,2560) : 0
(0,2240):(518,2560) : 0
ADDHX4
--pins(6)
S
use :  
dir : o
shape : 
(5484,316):(5648,478) : 0
(4314,316):(5484,426) : 0
(3036,1422):(5432,1530) : 0
(4192,316):(4314,784) : 0
(4086,600):(4192,784) : 0
(3076,674):(4086,784) : 0
(3036,600):(3076,1266) : 0
(2914,600):(3036,1530) : 0
(2874,600):(2914,1266) : 0
(2534,1422):(2914,1530) : 0
(2768,626):(2874,810) : 0
CO
use :  
dir : o
shape : 
(9296,1134):(9376,1800) : 0
(9174,676):(9296,1800) : 0
(9074,676):(9174,786) : 0
(8832,1330):(9174,1440) : 0
B
use :  
dir : i
shape : 
(4476,926):(5280,1036) : 0
(4468,926):(4476,1236) : 0
(4346,926):(4468,1254) : 0
(4314,1126):(4346,1254) : 0
(3388,1126):(4314,1236) : 0
A
use :  
dir : i
shape : 
(6576,976):(8222,1086) : 0
(6454,878):(6576,1086) : 0
(6414,878):(6454,988) : 0
VSS
use : g
dir : b
shape : 
(9594,-160):(9800,160) : 0
(9412,-160):(9594,428) : 0
(8914,-160):(9412,160) : 0
(8734,-160):(8914,428) : 0
(8202,-160):(8734,160) : 0
(8020,-160):(8202,422) : 0
(7522,-160):(8020,160) : 0
(7342,-160):(7522,422) : 0
(6844,-160):(7342,160) : 0
(6664,-160):(6844,396) : 0
(2482,-160):(6664,160) : 0
(2302,-160):(2482,244) : 0
(1654,-160):(2302,160) : 0
(1474,-160):(1654,244) : 0
(954,-160):(1474,160) : 0
(774,-160):(954,428) : 0
(276,-160):(774,160) : 0
(96,-160):(276,422) : 0
(0,-160):(96,160) : 0
VDD
use : p
dir : b
shape : 
(9410,2240):(9800,2560) : 0
(9172,2156):(9410,2560) : 0
(8662,2240):(9172,2560) : 0
(8482,1978):(8662,2560) : 0
(7970,2240):(8482,2560) : 0
(7790,1978):(7970,2560) : 0
(7292,2240):(7790,2560) : 0
(7112,1978):(7292,2560) : 0
(6590,2240):(7112,2560) : 0
(6408,2156):(6590,2560) : 0
(5762,2240):(6408,2560) : 0
(5582,2156):(5762,2560) : 0
(2376,2240):(5582,2560) : 0
(2196,2156):(2376,2560) : 0
(1654,2240):(2196,2560) : 0
(1474,2156):(1654,2560) : 0
(954,2240):(1474,2560) : 0
(774,1978):(954,2560) : 0
(276,2240):(774,2560) : 0
(96,1978):(276,2560) : 0
(0,2240):(96,2560) : 0
ADDHX2
--pins(6)
S
use :  
dir : o
shape : 
(3078,612):(3202,784) : 0
(2284,1348):(3156,1510) : 0
(1894,638):(3078,748) : 0
(2018,1374):(2284,1510) : 0
(1758,1374):(2018,1522) : 0
(1788,612):(1894,748) : 0
(1758,612):(1788,774) : 0
(1636,612):(1758,1522) : 0
(1606,612):(1636,774) : 0
(1624,1338):(1636,1522) : 0
CO
use :  
dir : o
shape : 
(5970,648):(6198,810) : 0
(5928,648):(5970,878) : 0
(5934,1252):(5964,1466) : 0
(5928,1252):(5934,1522) : 0
(5804,700):(5928,1522) : 0
(5780,1252):(5804,1466) : 0
B
use :  
dir : i
shape : 
(2772,876):(2954,1038) : 0
(2728,876):(2772,1012) : 0
(2604,878):(2728,1012) : 0
(2208,902):(2604,1012) : 0
(2084,902):(2208,1238) : 0
(2026,1076):(2084,1238) : 0
A
use :  
dir : i
shape : 
(4506,908):(5050,1070) : 0
(4382,878):(4506,1070) : 0
(4108,908):(4382,1070) : 0
VSS
use : g
dir : b
shape : 
(5810,-160):(6400,160) : 0
(5626,-160):(5810,422) : 0
(5132,-160):(5626,160) : 0
(4948,-160):(5132,440) : 0
(4442,-160):(4948,160) : 0
(4258,-160):(4442,440) : 0
(992,-160):(4258,160) : 0
(808,-160):(992,244) : 0
(280,-160):(808,160) : 0
(96,-160):(280,430) : 0
(0,-160):(96,160) : 0
VDD
use : p
dir : b
shape : 
(5618,2240):(6400,2560) : 0
(5436,1978):(5618,2560) : 0
(4896,2240):(5436,2560) : 0
(4714,1978):(4896,2560) : 0
(4208,2240):(4714,2560) : 0
(4024,2004):(4208,2560) : 0
(3534,2240):(4024,2560) : 0
(3350,2130):(3534,2560) : 0
(992,2240):(3350,2560) : 0
(808,2156):(992,2560) : 0
(280,2240):(808,2560) : 0
(96,2004):(280,2560) : 0
(0,2240):(96,2560) : 0
ADDHX1
--pins(6)
S
use :  
dir : o
shape : 
(2124,634):(2246,1534) : 0
(1904,634):(2124,742) : 0
(1720,1352):(2124,1534) : 0
(1782,576):(1904,742) : 0
(1598,1352):(1720,1776) : 0
CO
use :  
dir : o
shape : 
(4036,878):(4086,988) : 0
(3924,658):(4036,988) : 0
(3914,658):(3924,1484) : 0
(3802,878):(3914,1484) : 0
(3726,1374):(3802,1484) : 0
(3604,1374):(3726,1890) : 0
B
use :  
dir : i
shape : 
(3094,1200):(3216,1640) : 0
(2736,1530):(3094,1640) : 0
(2614,1530):(2736,2016) : 0
(1476,1908):(2614,2016) : 0
(1880,858):(2002,1200) : 0
(1476,1090):(1880,1200) : 0
(1354,1090):(1476,2016) : 0
(1164,1090):(1354,1266) : 0
(1122,1090):(1164,1226) : 0
(942,1064):(1122,1226) : 0
A
use :  
dir : i
shape : 
(2368,866):(2692,1066) : 0
VSS
use : g
dir : b
shape : 
(3792,-160):(4200,160) : 0
(3670,-160):(3792,666) : 0
(2718,-160):(3670,160) : 0
(3614,566):(3670,666) : 0
(3492,566):(3614,790) : 0
(2538,-160):(2718,244) : 0
(722,-160):(2538,160) : 0
(540,-160):(722,244) : 0
(0,-160):(540,160) : 0
VDD
use : p
dir : b
shape : 
(3436,2240):(4200,2560) : 0
(3256,2156):(3436,2560) : 0
(2534,2240):(3256,2560) : 0
(2354,2156):(2534,2560) : 0
(678,2240):(2354,2560) : 0
(498,2156):(678,2560) : 0
(0,2240):(498,2560) : 0
ADDFX2
--pins(7)
S
use :  
dir : o
shape : 
(7114,612):(7138,848) : 0
(7114,1330):(7130,1492) : 0
(6992,612):(7114,1492) : 0
(6956,612):(6992,848) : 0
(6948,1330):(6992,1492) : 0
(6810,612):(6956,722) : 0
CO
use :  
dir : o
shape : 
(6278,680):(6410,842) : 0
(6278,1330):(6398,1492) : 0
(6156,680):(6278,1492) : 0
(6106,1146):(6156,1254) : 0
CI
use :  
dir : i
shape : 
(4922,866):(5064,976) : 0
(4800,866):(4922,1534) : 0
(4592,1364):(4800,1534) : 0
B
use :  
dir : i
shape : 
(238,972):(406,1134) : 0
(224,972):(238,1254) : 0
(114,1024):(224,1254) : 0
A
use :  
dir : i
shape : 
(2080,1120):(2582,1280) : 0
VSS
use : g
dir : b
shape : 
(6776,-160):(7400,160) : 0
(6594,-160):(6776,244) : 0
(5382,-160):(6594,160) : 0
(5200,-160):(5382,244) : 0
(2522,-160):(5200,160) : 0
(2342,-160):(2522,398) : 0
(686,-160):(2342,160) : 0
(504,-160):(686,244) : 0
(0,-160):(504,160) : 0
VDD
use : p
dir : b
shape : 
(6768,2240):(7400,2560) : 0
(6586,2156):(6768,2560) : 0
(4770,2240):(6586,2560) : 0
(4588,2156):(4770,2560) : 0
(640,2240):(4588,2560) : 0
(460,2156):(640,2560) : 0
(0,2240):(460,2560) : 0
ADDFX1
--pins(7)
S
use :  
dir : o
shape : 
(7246,612):(7286,722) : 0
(7186,612):(7246,878) : 0
(7186,1254):(7246,1716) : 0
(7064,612):(7186,1716) : 0
CO
use :  
dir : o
shape : 
(6410,1134):(6580,1266) : 0
(6398,680):(6410,1266) : 0
(6276,680):(6398,1492) : 0
(6228,680):(6276,842) : 0
(6218,1330):(6276,1492) : 0
CI
use :  
dir : i
shape : 
(4922,866):(5064,976) : 0
(4800,866):(4922,1534) : 0
(4592,1364):(4800,1534) : 0
B
use :  
dir : i
shape : 
(238,972):(406,1134) : 0
(224,972):(238,1254) : 0
(114,1024):(224,1254) : 0
A
use :  
dir : i
shape : 
(2080,1120):(2582,1280) : 0
VSS
use : g
dir : b
shape : 
(6818,-160):(7400,160) : 0
(6636,-160):(6818,740) : 0
(5382,-160):(6636,160) : 0
(5200,-160):(5382,244) : 0
(2522,-160):(5200,160) : 0
(2342,-160):(2522,398) : 0
(686,-160):(2342,160) : 0
(504,-160):(686,244) : 0
(0,-160):(504,160) : 0
VDD
use : p
dir : b
shape : 
(6820,2240):(7400,2560) : 0
(6640,1902):(6820,2560) : 0
(4770,2240):(6640,2560) : 0
(4588,2156):(4770,2560) : 0
(640,2240):(4588,2560) : 0
(460,2156):(640,2560) : 0
(0,2240):(460,2560) : 0
ADDFHX4
--pins(7)
S
use :  
dir : o
shape : 
(11698,866):(11778,1534) : 0
(11576,666):(11698,1534) : 0
(11466,666):(11576,828) : 0
(11466,1342):(11576,1504) : 0
CO
use :  
dir : o
shape : 
(11002,866):(11080,1534) : 0
(10880,692):(11002,1534) : 0
(10790,692):(10880,802) : 0
(10788,1342):(10880,1504) : 0
CI
use :  
dir : i
shape : 
(10032,1134):(10384,1316) : 0
B
use :  
dir : i
shape : 
(7206,1270):(7430,1430) : 0
(7084,1270):(7206,1522) : 0
(6754,1270):(7084,1430) : 0
A
use :  
dir : i
shape : 
(382,866):(658,1142) : 0
VSS
use : g
dir : b
shape : 
(11984,-160):(12200,160) : 0
(11804,-160):(11984,466) : 0
(11308,-160):(11804,160) : 0
(11128,-160):(11308,466) : 0
(10590,-160):(11128,160) : 0
(10410,-160):(10590,244) : 0
(7172,-160):(10410,160) : 0
(6992,-160):(7172,244) : 0
(1728,-160):(6992,160) : 0
(1548,-160):(1728,244) : 0
(660,-160):(1548,160) : 0
(480,-160):(660,244) : 0
(0,-160):(480,160) : 0
VDD
use : p
dir : b
shape : 
(11986,2240):(12200,2560) : 0
(11806,1976):(11986,2560) : 0
(11308,2240):(11806,2560) : 0
(11128,1976):(11308,2560) : 0
(10628,2240):(11128,2560) : 0
(10450,1978):(10628,2560) : 0
(9936,2240):(10450,2560) : 0
(9700,2156):(9936,2560) : 0
(7442,2240):(9700,2560) : 0
(7262,1940):(7442,2560) : 0
(6680,2240):(7262,2560) : 0
(6502,1940):(6680,2560) : 0
(1932,2240):(6502,2560) : 0
(1754,1822):(1932,2560) : 0
(764,2240):(1754,2560) : 0
(584,1934):(764,2560) : 0
(0,2240):(584,2560) : 0
ADDFHX2
--pins(7)
S
use :  
dir : o
shape : 
(11594,438):(11690,988) : 0
(11594,1254):(11624,1916) : 0
(11510,438):(11594,1916) : 0
(11474,714):(11510,1916) : 0
(11446,1308):(11474,1916) : 0
CO
use :  
dir : o
shape : 
(10932,662):(11028,824) : 0
(10848,662):(10932,1522) : 0
(10812,688):(10848,1522) : 0
(10524,1412):(10812,1522) : 0
CI
use :  
dir : i
shape : 
(9988,1092):(10338,1298) : 0
B
use :  
dir : i
shape : 
(7176,1270):(7398,1430) : 0
(7054,1270):(7176,1522) : 0
(6726,1270):(7054,1430) : 0
A
use :  
dir : i
shape : 
(382,866):(654,1142) : 0
VSS
use : g
dir : b
shape : 
(11310,-160):(11800,160) : 0
(11132,-160):(11310,422) : 0
(10628,-160):(11132,160) : 0
(10448,-160):(10628,244) : 0
(7140,-160):(10448,160) : 0
(6962,-160):(7140,244) : 0
(1762,-160):(6962,160) : 0
(1582,-160):(1762,244) : 0
(700,-160):(1582,160) : 0
(520,-160):(700,244) : 0
(0,-160):(520,160) : 0
VDD
use : p
dir : b
shape : 
(11246,2240):(11800,2560) : 0
(11066,1976):(11246,2560) : 0
(10582,2240):(11066,2560) : 0
(10404,1976):(10582,2560) : 0
(9880,2240):(10404,2560) : 0
(9668,2156):(9880,2560) : 0
(7410,2240):(9668,2560) : 0
(7230,1940):(7410,2560) : 0
(6652,2240):(7230,2560) : 0
(6474,1940):(6652,2560) : 0
(1924,2240):(6474,2560) : 0
(1746,1822):(1924,2560) : 0
(760,2240):(1746,2560) : 0
(582,1934):(760,2560) : 0
(0,2240):(582,2560) : 0
ADDFHX1
--pins(7)
S
use :  
dir : o
shape : 
(7876,878):(7886,988) : 0
(7754,652):(7876,1676) : 0
CO
use :  
dir : o
shape : 
(7180,878):(7192,988) : 0
(7060,652):(7180,1754) : 0
(6910,1646):(7060,1754) : 0
CI
use :  
dir : i
shape : 
(6650,1400):(6844,1522) : 0
(6530,1120):(6650,1522) : 0
B
use :  
dir : i
shape : 
(3638,1400):(4060,1608) : 0
A
use :  
dir : i
shape : 
(376,878):(582,1186) : 0
VSS
use : g
dir : b
shape : 
(7610,-160):(8000,160) : 0
(7430,-160):(7610,244) : 0
(6896,-160):(7430,160) : 0
(6716,-160):(6896,244) : 0
(4034,-160):(6716,160) : 0
(3856,-160):(4034,244) : 0
(928,-160):(3856,160) : 0
(748,-160):(928,244) : 0
(0,-160):(748,160) : 0
VDD
use : p
dir : b
shape : 
(7488,2240):(8000,2560) : 0
(7310,2156):(7488,2560) : 0
(6314,2240):(7310,2560) : 0
(6134,2156):(6314,2560) : 0
(3944,2240):(6134,2560) : 0
(3766,1966):(3944,2560) : 0
(1256,2240):(3766,2560) : 0
(1078,1788):(1256,2560) : 0
(654,2240):(1078,2560) : 0
(474,1818):(654,2560) : 0
(0,2240):(474,2560) : 0
XOR3X4
--pins(6)
Y
use :  
dir : o
shape : 
(9954,1400):(9980,2066) : 0
(9928,454):(9954,2066) : 0
(9832,398):(9928,2066) : 0
(9748,398):(9832,784) : 0
(9780,1304):(9832,2066) : 0
(9770,1304):(9780,1466) : 0
C
use :  
dir : i
shape : 
(9114,1872):(9292,2034) : 0
(8900,1924):(9114,2034) : 0
(8780,1924):(8900,2054) : 0
B
use :  
dir : i
shape : 
(6304,1274):(6360,1436) : 0
(6182,750):(6304,1436) : 0
(6050,750):(6182,1000) : 0
(6006,878):(6050,1000) : 0
A
use :  
dir : i
shape : 
(580,1052):(772,1214) : 0
(460,1052):(580,1254) : 0
(346,1052):(460,1214) : 0
VSS
use : g
dir : b
shape : 
(10306,-160):(10400,160) : 0
(10126,-160):(10306,754) : 0
(9528,-160):(10126,160) : 0
(9350,-160):(9528,270) : 0
(4924,-160):(9350,160) : 0
(4746,-160):(4924,244) : 0
(4020,-160):(4746,160) : 0
(3842,-160):(4020,244) : 0
(3202,-160):(3842,160) : 0
(3022,-160):(3202,244) : 0
(672,-160):(3022,160) : 0
(494,-160):(672,718) : 0
(0,-160):(494,160) : 0
VDD
use : p
dir : b
shape : 
(10306,2240):(10400,2560) : 0
(10126,1906):(10306,2560) : 0
(9592,2240):(10126,2560) : 0
(9412,1906):(9592,2560) : 0
(4730,2240):(9412,2560) : 0
(4552,2130):(4730,2560) : 0
(3932,2240):(4552,2560) : 0
(3752,2042):(3932,2560) : 0
(3134,2240):(3752,2560) : 0
(2954,2042):(3134,2560) : 0
(662,2240):(2954,2560) : 0
(484,1906):(662,2560) : 0
(0,2240):(484,2560) : 0
XOR3X2
--pins(6)
Y
use :  
dir : o
shape : 
(6304,454):(6330,1440) : 0
(6284,398):(6304,1466) : 0
(6206,398):(6284,1522) : 0
(6120,398):(6206,784) : 0
(6160,1304):(6206,1522) : 0
(6120,1304):(6160,1466) : 0
C
use :  
dir : i
shape : 
(5344,1576):(5630,1800) : 0
B
use :  
dir : i
shape : 
(3784,1146):(3796,1254) : 0
(3726,1146):(3784,1538) : 0
(3602,852):(3726,1538) : 0
(3428,852):(3602,1014) : 0
A
use :  
dir : i
shape : 
(240,1052):(442,1214) : 0
(116,1052):(240,1254) : 0
(76,1052):(116,1214) : 0
VSS
use : g
dir : b
shape : 
(5894,-160):(6400,160) : 0
(5710,-160):(5894,270) : 0
(1990,-160):(5710,160) : 0
(1808,-160):(1990,358) : 0
(280,-160):(1808,160) : 0
(96,-160):(280,718) : 0
(0,-160):(96,160) : 0
VDD
use : p
dir : b
shape : 
(5936,2240):(6400,2560) : 0
(5754,1906):(5936,2560) : 0
(1904,2240):(5754,2560) : 0
(1722,2022):(1904,2560) : 0
(324,2240):(1722,2560) : 0
(140,1906):(324,2560) : 0
(0,2240):(140,2560) : 0
XNOR3X4
--pins(6)
Y
use :  
dir : o
shape : 
(9954,1400):(9980,2066) : 0
(9928,454):(9954,2066) : 0
(9832,398):(9928,2066) : 0
(9748,398):(9832,784) : 0
(9780,1304):(9832,2066) : 0
(9770,1304):(9780,1466) : 0
C
use :  
dir : i
shape : 
(9114,1872):(9292,2034) : 0
(8900,1924):(9114,2034) : 0
(8780,1924):(8900,2054) : 0
B
use :  
dir : i
shape : 
(6282,1274):(6340,1436) : 0
(6162,750):(6282,1436) : 0
(6050,750):(6162,1000) : 0
(6006,878):(6050,1000) : 0
A
use :  
dir : i
shape : 
(580,1052):(772,1214) : 0
(460,1052):(580,1254) : 0
(346,1052):(460,1214) : 0
VSS
use : g
dir : b
shape : 
(10306,-160):(10400,160) : 0
(10126,-160):(10306,754) : 0
(9528,-160):(10126,160) : 0
(9350,-160):(9528,270) : 0
(4924,-160):(9350,160) : 0
(4746,-160):(4924,244) : 0
(4020,-160):(4746,160) : 0
(3842,-160):(4020,244) : 0
(3202,-160):(3842,160) : 0
(3022,-160):(3202,244) : 0
(672,-160):(3022,160) : 0
(494,-160):(672,718) : 0
(0,-160):(494,160) : 0
VDD
use : p
dir : b
shape : 
(10306,2240):(10400,2560) : 0
(10126,1906):(10306,2560) : 0
(9592,2240):(10126,2560) : 0
(9412,1906):(9592,2560) : 0
(4730,2240):(9412,2560) : 0
(4552,2130):(4730,2560) : 0
(3932,2240):(4552,2560) : 0
(3752,2042):(3932,2560) : 0
(3134,2240):(3752,2560) : 0
(2954,2042):(3134,2560) : 0
(662,2240):(2954,2560) : 0
(484,1906):(662,2560) : 0
(0,2240):(484,2560) : 0
XNOR3X2
--pins(6)
Y
use :  
dir : o
shape : 
(6304,454):(6330,1440) : 0
(6284,398):(6304,1466) : 0
(6206,398):(6284,1522) : 0
(6120,398):(6206,784) : 0
(6160,1304):(6206,1522) : 0
(6120,1304):(6160,1466) : 0
C
use : 
dir : i
shape : 
(5344,1576):(5630,1800) : 0
B
use : �
dir : i
shape : 
(3784,1146):(3796,1254) : 0
(3726,1146):(3784,1538) : 0
(3602,852):(3726,1538) : 0
(3428,852):(3602,1014) : 0
A
use : 
dir : i
shape : 
(240,1052):(442,1214) : 0
(116,1052):(240,1254) : 0
(76,1052):(116,1214) : 0
VSS
use : g
dir : b
shape : 
(5894,-160):(6400,160) : 0
(5710,-160):(5894,270) : 0
(1990,-160):(5710,160) : 0
(1808,-160):(1990,358) : 0
(280,-160):(1808,160) : 0
(96,-160):(280,718) : 0
(0,-160):(96,160) : 0
VDD
use : p
dir : b
shape : 
(5936,2240):(6400,2560) : 0
(5754,1906):(5936,2560) : 0
(1904,2240):(5754,2560) : 0
(1722,2022):(1904,2560) : 0
(324,2240):(1722,2560) : 0
(140,1906):(324,2560) : 0
(0,2240):(140,2560) : 0
ram_256x16A
--pins(46)
A[0]
use : s
dir : i
shape : 
(61996,3440):(62216,3860) : 0
(61996,3440):(62216,3860) : 1
(61996,3440):(62216,3860) : 2
(61996,3440):(62216,3860) : 3
A[1]
use : s
dir : i
shape : 
(61264,3440):(61484,3860) : 0
(61264,3440):(61484,3860) : 1
(61264,3440):(61484,3860) : 2
(61264,3440):(61484,3860) : 3
A[2]
use : s
dir : i
shape : 
(60236,3440):(60456,3860) : 0
(60236,3440):(60456,3860) : 1
(60236,3440):(60456,3860) : 2
(60236,3440):(60456,3860) : 3
A[3]
use : s
dir : i
shape : 
(59504,3440):(59724,3860) : 0
(59504,3440):(59724,3860) : 1
(59504,3440):(59724,3860) : 2
(59504,3440):(59724,3860) : 3
A[4]
use : s
dir : i
shape : 
(57744,3440):(57964,3860) : 0
(57744,3440):(57964,3860) : 1
(57744,3440):(57964,3860) : 2
(57744,3440):(57964,3860) : 3
A[5]
use : s
dir : i
shape : 
(56716,3440):(56936,3860) : 0
(56716,3440):(56936,3860) : 1
(56716,3440):(56936,3860) : 2
(56716,3440):(56936,3860) : 3
A[6]
use : s
dir : i
shape : 
(55984,3440):(56204,3860) : 0
(55984,3440):(56204,3860) : 1
(55984,3440):(56204,3860) : 2
(55984,3440):(56204,3860) : 3
A[7]
use : s
dir : i
shape : 
(54224,3440):(54444,3860) : 0
(54224,3440):(54444,3860) : 1
(54224,3440):(54444,3860) : 2
(54224,3440):(54444,3860) : 3
CEN
use : s
dir : i
shape : 
(63736,3440):(63956,3860) : 0
(63736,3440):(63956,3860) : 1
(63736,3440):(63956,3860) : 2
(63736,3440):(63956,3860) : 3
CLK
use : c
dir : i
shape : 
(66642,3440):(66862,3860) : 0
(66642,3440):(66862,3860) : 1
(66642,3440):(66862,3860) : 2
(66642,3440):(66862,3860) : 3
D[0]
use : s
dir : i
shape : 
(9092,3440):(9312,3860) : 0
(9092,3440):(9312,3860) : 1
(9092,3440):(9312,3860) : 2
(9092,3440):(9312,3860) : 3
D[10]
use : s
dir : i
shape : 
(83896,3440):(84116,3860) : 0
(83896,3440):(84116,3860) : 1
(83896,3440):(84116,3860) : 2
(83896,3440):(84116,3860) : 3
D[11]
use : s
dir : i
shape : 
(86060,3440):(86280,3860) : 0
(86060,3440):(86280,3860) : 1
(86060,3440):(86280,3860) : 2
(86060,3440):(86280,3860) : 3
D[12]
use : s
dir : i
shape : 
(96032,3440):(96252,3860) : 0
(96032,3440):(96252,3860) : 1
(96032,3440):(96252,3860) : 2
(96032,3440):(96252,3860) : 3
D[13]
use : s
dir : i
shape : 
(98196,3440):(98416,3860) : 0
(98196,3440):(98416,3860) : 1
(98196,3440):(98416,3860) : 2
(98196,3440):(98416,3860) : 3
D[14]
use : s
dir : i
shape : 
(108168,3440):(108388,3860) : 0
(108168,3440):(108388,3860) : 1
(108168,3440):(108388,3860) : 2
(108168,3440):(108388,3860) : 3
D[15]
use : s
dir : i
shape : 
(110332,3440):(110552,3860) : 0
(110332,3440):(110552,3860) : 1
(110332,3440):(110552,3860) : 2
(110332,3440):(110552,3860) : 3
D[1]
use : s
dir : i
shape : 
(11256,3440):(11476,3860) : 0
(11256,3440):(11476,3860) : 1
(11256,3440):(11476,3860) : 2
(11256,3440):(11476,3860) : 3
D[2]
use : s
dir : i
shape : 
(21228,3440):(21448,3860) : 0
(21228,3440):(21448,3860) : 1
(21228,3440):(21448,3860) : 2
(21228,3440):(21448,3860) : 3
D[3]
use : s
dir : i
shape : 
(23392,3440):(23612,3860) : 0
(23392,3440):(23612,3860) : 1
(23392,3440):(23612,3860) : 2
(23392,3440):(23612,3860) : 3
D[4]
use : s
dir : i
shape : 
(33364,3440):(33584,3860) : 0
(33364,3440):(33584,3860) : 1
(33364,3440):(33584,3860) : 2
(33364,3440):(33584,3860) : 3
D[5]
use : s
dir : i
shape : 
(35528,3440):(35748,3860) : 0
(35528,3440):(35748,3860) : 1
(35528,3440):(35748,3860) : 2
(35528,3440):(35748,3860) : 3
D[6]
use : s
dir : i
shape : 
(45500,3440):(45720,3860) : 0
(45500,3440):(45720,3860) : 1
(45500,3440):(45720,3860) : 2
(45500,3440):(45720,3860) : 3
D[7]
use : s
dir : i
shape : 
(47664,3440):(47884,3860) : 0
(47664,3440):(47884,3860) : 1
(47664,3440):(47884,3860) : 2
(47664,3440):(47884,3860) : 3
D[8]
use : s
dir : i
shape : 
(71760,3440):(71980,3860) : 0
(71760,3440):(71980,3860) : 1
(71760,3440):(71980,3860) : 2
(71760,3440):(71980,3860) : 3
D[9]
use : s
dir : i
shape : 
(73924,3440):(74144,3860) : 0
(73924,3440):(74144,3860) : 1
(73924,3440):(74144,3860) : 2
(73924,3440):(74144,3860) : 3
OEN
use : s
dir : i
shape : 
(66040,3440):(66260,3860) : 0
(66040,3440):(66260,3860) : 1
(66040,3440):(66260,3860) : 2
(66040,3440):(66260,3860) : 3
Q[0]
use : s
dir :  
shape : 
(7996,3440):(8216,3860) : 0
(7996,3440):(8216,3860) : 1
(7996,3440):(8216,3860) : 2
(7996,3440):(8216,3860) : 3
Q[10]
use : s
dir :  
shape : 
(82840,3440):(83060,3860) : 0
(82840,3440):(83060,3860) : 1
(82840,3440):(83060,3860) : 2
(82840,3440):(83060,3860) : 3
Q[11]
use : s
dir :  
shape : 
(87116,3440):(87336,3860) : 0
(87116,3440):(87336,3860) : 1
(87116,3440):(87336,3860) : 2
(87116,3440):(87336,3860) : 3
Q[12]
use : s
dir :  
shape : 
(94976,3440):(95196,3860) : 0
(94976,3440):(95196,3860) : 1
(94976,3440):(95196,3860) : 2
(94976,3440):(95196,3860) : 3
Q[13]
use : s
dir :  
shape : 
(99252,3440):(99472,3860) : 0
(99252,3440):(99472,3860) : 1
(99252,3440):(99472,3860) : 2
(99252,3440):(99472,3860) : 3
Q[14]
use : s
dir :  
shape : 
(107112,3440):(107332,3860) : 0
(107112,3440):(107332,3860) : 1
(107112,3440):(107332,3860) : 2
(107112,3440):(107332,3860) : 3
Q[15]
use : s
dir :  
shape : 
(111408,3440):(111628,3860) : 0
(111408,3440):(111628,3860) : 1
(111408,3440):(111628,3860) : 2
(111408,3440):(111628,3860) : 3
Q[1]
use : s
dir :  
shape : 
(12312,3440):(12532,3860) : 0
(12312,3440):(12532,3860) : 1
(12312,3440):(12532,3860) : 2
(12312,3440):(12532,3860) : 3
Q[2]
use : s
dir :  
shape : 
(20172,3440):(20392,3860) : 0
(20172,3440):(20392,3860) : 1
(20172,3440):(20392,3860) : 2
(20172,3440):(20392,3860) : 3
Q[3]
use : s
dir :  
shape : 
(24448,3440):(24668,3860) : 0
(24448,3440):(24668,3860) : 1
(24448,3440):(24668,3860) : 2
(24448,3440):(24668,3860) : 3
Q[4]
use : s
dir :  
shape : 
(32308,3440):(32528,3860) : 0
(32308,3440):(32528,3860) : 1
(32308,3440):(32528,3860) : 2
(32308,3440):(32528,3860) : 3
Q[5]
use : s
dir :  
shape : 
(36584,3440):(36804,3860) : 0
(36584,3440):(36804,3860) : 1
(36584,3440):(36804,3860) : 2
(36584,3440):(36804,3860) : 3
Q[6]
use : s
dir :  
shape : 
(44444,3440):(44664,3860) : 0
(44444,3440):(44664,3860) : 1
(44444,3440):(44664,3860) : 2
(44444,3440):(44664,3860) : 3
Q[7]
use : s
dir :  
shape : 
(48720,3440):(48940,3860) : 0
(48720,3440):(48940,3860) : 1
(48720,3440):(48940,3860) : 2
(48720,3440):(48940,3860) : 3
Q[8]
use : s
dir :  
shape : 
(70704,3440):(70924,3860) : 0
(70704,3440):(70924,3860) : 1
(70704,3440):(70924,3860) : 2
(70704,3440):(70924,3860) : 3
Q[9]
use : s
dir :  
shape : 
(74980,3440):(75200,3860) : 0
(74980,3440):(75200,3860) : 1
(74980,3440):(75200,3860) : 2
(74980,3440):(75200,3860) : 3
WEN
use : s
dir : i
shape : 
(64312,3440):(64532,3860) : 0
(64312,3440):(64532,3860) : 1
(64312,3440):(64532,3860) : 2
(64312,3440):(64532,3860) : 3
VDD
use : p
dir : b
shape : 
(0,36448):(119644,37848) : 4
(0,0):(119644,1400) : 4
(118244,0):(119644,37848) : 3
(0,0):(1400,37848) : 3
VSS
use : g
dir : b
shape : 
(1720,34728):(117924,36128) : 4
(1720,1720):(117924,3120) : 4
(116524,1720):(117924,36128) : 3
(1720,1720):(3120,36128) : 3
rom_512x16A
--pins(29)
A[0]
use : s
dir : i
shape : 
(17740,4240):(17962,4660) : 0
(17740,4240):(17962,4660) : 1
(17740,4240):(17962,4660) : 2
(17740,4240):(17962,4660) : 3
A[1]
use : s
dir : i
shape : 
(16842,4240):(17062,4660) : 0
(16842,4240):(17062,4660) : 1
(16842,4240):(17062,4660) : 2
(16842,4240):(17062,4660) : 3
A[2]
use : s
dir : i
shape : 
(15942,4240):(16162,4660) : 0
(15942,4240):(16162,4660) : 1
(15942,4240):(16162,4660) : 2
(15942,4240):(16162,4660) : 3
A[3]
use : s
dir : i
shape : 
(14142,4240):(14362,4660) : 0
(14142,4240):(14362,4660) : 1
(14142,4240):(14362,4660) : 2
(14142,4240):(14362,4660) : 3
A[4]
use : s
dir : i
shape : 
(12342,4240):(12562,4660) : 0
(12342,4240):(12562,4660) : 1
(12342,4240):(12562,4660) : 2
(12342,4240):(12562,4660) : 3
A[5]
use : s
dir : i
shape : 
(11442,4240):(11662,4660) : 0
(11442,4240):(11662,4660) : 1
(11442,4240):(11662,4660) : 2
(11442,4240):(11662,4660) : 3
A[6]
use : s
dir : i
shape : 
(10542,4240):(10762,4660) : 0
(10542,4240):(10762,4660) : 1
(10542,4240):(10762,4660) : 2
(10542,4240):(10762,4660) : 3
A[7]
use : s
dir : i
shape : 
(8740,4240):(8962,4660) : 0
(8740,4240):(8962,4660) : 1
(8740,4240):(8962,4660) : 2
(8740,4240):(8962,4660) : 3
A[8]
use : s
dir : i
shape : 
(7842,4240):(8060,4660) : 0
(7842,4240):(8060,4660) : 1
(7842,4240):(8060,4660) : 2
(7842,4240):(8060,4660) : 3
CEN
use : s
dir : i
shape : 
(22404,4240):(22624,4660) : 0
(22404,4240):(22624,4660) : 1
(22404,4240):(22624,4660) : 2
(22404,4240):(22624,4660) : 3
CLK
use : c
dir : i
shape : 
(22064,4240):(22284,4660) : 0
(22064,4240):(22284,4660) : 1
(22064,4240):(22284,4660) : 2
(22064,4240):(22284,4660) : 3
Q[0]
use : s
dir :  
shape : 
(28314,4240):(28536,4660) : 0
(28314,4240):(28536,4660) : 1
(28314,4240):(28536,4660) : 2
(28314,4240):(28536,4660) : 3
Q[10]
use : s
dir :  
shape : 
(55096,4240):(55314,4660) : 0
(55096,4240):(55314,4660) : 1
(55096,4240):(55314,4660) : 2
(55096,4240):(55314,4660) : 3
Q[11]
use : s
dir :  
shape : 
(55708,4240):(55926,4660) : 0
(55708,4240):(55926,4660) : 1
(55708,4240):(55926,4660) : 2
(55708,4240):(55926,4660) : 3
Q[12]
use : s
dir :  
shape : 
(60452,4240):(60672,4660) : 0
(60452,4240):(60672,4660) : 1
(60452,4240):(60672,4660) : 2
(60452,4240):(60672,4660) : 3
Q[13]
use : s
dir :  
shape : 
(61064,4240):(61284,4660) : 0
(61064,4240):(61284,4660) : 1
(61064,4240):(61284,4660) : 2
(61064,4240):(61284,4660) : 3
Q[14]
use : s
dir :  
shape : 
(65808,4240):(66028,4660) : 0
(65808,4240):(66028,4660) : 1
(65808,4240):(66028,4660) : 2
(65808,4240):(66028,4660) : 3
Q[15]
use : s
dir :  
shape : 
(66420,4240):(66640,4660) : 0
(66420,4240):(66640,4660) : 1
(66420,4240):(66640,4660) : 2
(66420,4240):(66640,4660) : 3
Q[1]
use : s
dir :  
shape : 
(28926,4240):(29148,4660) : 0
(28926,4240):(29148,4660) : 1
(28926,4240):(29148,4660) : 2
(28926,4240):(29148,4660) : 3
Q[2]
use : s
dir :  
shape : 
(33670,4240):(33892,4660) : 0
(33670,4240):(33892,4660) : 1
(33670,4240):(33892,4660) : 2
(33670,4240):(33892,4660) : 3
Q[3]
use : s
dir :  
shape : 
(34284,4240):(34504,4660) : 0
(34284,4240):(34504,4660) : 1
(34284,4240):(34504,4660) : 2
(34284,4240):(34504,4660) : 3
Q[4]
use : s
dir :  
shape : 
(39028,4240):(39248,4660) : 0
(39028,4240):(39248,4660) : 1
(39028,4240):(39248,4660) : 2
(39028,4240):(39248,4660) : 3
Q[5]
use : s
dir :  
shape : 
(39640,4240):(39860,4660) : 0
(39640,4240):(39860,4660) : 1
(39640,4240):(39860,4660) : 2
(39640,4240):(39860,4660) : 3
Q[6]
use : s
dir :  
shape : 
(44384,4240):(44604,4660) : 0
(44384,4240):(44604,4660) : 1
(44384,4240):(44604,4660) : 2
(44384,4240):(44604,4660) : 3
Q[7]
use : s
dir :  
shape : 
(44996,4240):(45216,4660) : 0
(44996,4240):(45216,4660) : 1
(44996,4240):(45216,4660) : 2
(44996,4240):(45216,4660) : 3
Q[8]
use : s
dir :  
shape : 
(49740,4240):(49960,4660) : 0
(49740,4240):(49960,4660) : 1
(49740,4240):(49960,4660) : 2
(49740,4240):(49960,4660) : 3
Q[9]
use : s
dir :  
shape : 
(50350,4240):(50570,4660) : 0
(50350,4240):(50570,4660) : 1
(50350,4240):(50570,4660) : 2
(50350,4240):(50570,4660) : 3
VDD
use : p
dir : o
shape : 
(0,35568):(73634,37368) : 4
(0,0):(73634,1800) : 4
(71834,0):(73634,37368) : 3
(0,0):(1800,37368) : 3
VSS
use : g
dir : o
shape : 
(2120,33450):(71514,35250) : 4
(2120,2120):(71514,3920) : 4
(69714,2120):(71514,35250) : 3
(2120,2120):(3920,35250) : 3
pllclk
--pins(11)
refclk
use :  
dir : i
shape : 
(0,30000):(520,30400) : 1
(0,30000):(520,30400) : 2
clk1x
use :  
dir : o
shape : 
(0,10000):(520,10400) : 1
(0,10000):(520,10400) : 2
clk2x
use :  
dir : o
shape : 
(0,12000):(520,12400) : 1
(0,12000):(520,12400) : 2
ibias
use :  
dir : i
shape : 
(0,36080):(520,36380) : 1
(0,36080):(520,36380) : 2
reset
use :  
dir : i
shape : 
(0,37008):(520,37308) : 1
(0,37008):(520,37308) : 2
vcom
use :  
dir : o
shape : 
(0,34244):(520,34544) : 1
(0,34244):(520,34544) : 2
vcop
use :  
dir : o
shape : 
(0,35172):(520,35472) : 1
(0,35172):(520,35472) : 2
AVSS
use : g
dir : b
shape : 
(29480,35692):(30000,36692) : 2
AVDD
use : p
dir : b
shape : 
(29480,32370):(30000,33372) : 2
VSS
use : g
dir : b
shape : 
(29480,4274):(30000,5274) : 2
VDD
use : p
dir : b
shape : 
(29480,954):(30000,1954) : 2
ram_128x16A
--pins(45)
A[0]
use : s
dir : i
shape : 
(61116,3440):(61336,3860) : 0
(61116,3440):(61336,3860) : 1
(61116,3440):(61336,3860) : 2
(61116,3440):(61336,3860) : 3
A[1]
use : s
dir : i
shape : 
(60384,3440):(60604,3860) : 0
(60384,3440):(60604,3860) : 1
(60384,3440):(60604,3860) : 2
(60384,3440):(60604,3860) : 3
A[2]
use : s
dir : i
shape : 
(59356,3440):(59576,3860) : 0
(59356,3440):(59576,3860) : 1
(59356,3440):(59576,3860) : 2
(59356,3440):(59576,3860) : 3
A[3]
use : s
dir : i
shape : 
(58624,3440):(58844,3860) : 0
(58624,3440):(58844,3860) : 1
(58624,3440):(58844,3860) : 2
(58624,3440):(58844,3860) : 3
A[4]
use : s
dir : i
shape : 
(56864,3440):(57084,3860) : 0
(56864,3440):(57084,3860) : 1
(56864,3440):(57084,3860) : 2
(56864,3440):(57084,3860) : 3
A[5]
use : s
dir : i
shape : 
(55836,3440):(56056,3860) : 0
(55836,3440):(56056,3860) : 1
(55836,3440):(56056,3860) : 2
(55836,3440):(56056,3860) : 3
A[6]
use : s
dir : i
shape : 
(55104,3440):(55324,3860) : 0
(55104,3440):(55324,3860) : 1
(55104,3440):(55324,3860) : 2
(55104,3440):(55324,3860) : 3
CEN
use : s
dir : i
shape : 
(62856,3440):(63076,3860) : 0
(62856,3440):(63076,3860) : 1
(62856,3440):(63076,3860) : 2
(62856,3440):(63076,3860) : 3
CLK
use : c
dir : i
shape : 
(65762,3440):(65982,3860) : 0
(65762,3440):(65982,3860) : 1
(65762,3440):(65982,3860) : 2
(65762,3440):(65982,3860) : 3
D[0]
use : s
dir : i
shape : 
(9092,3440):(9312,3860) : 0
(9092,3440):(9312,3860) : 1
(9092,3440):(9312,3860) : 2
(9092,3440):(9312,3860) : 3
D[10]
use : s
dir : i
shape : 
(83016,3440):(83236,3860) : 0
(83016,3440):(83236,3860) : 1
(83016,3440):(83236,3860) : 2
(83016,3440):(83236,3860) : 3
D[11]
use : s
dir : i
shape : 
(85180,3440):(85400,3860) : 0
(85180,3440):(85400,3860) : 1
(85180,3440):(85400,3860) : 2
(85180,3440):(85400,3860) : 3
D[12]
use : s
dir : i
shape : 
(95152,3440):(95372,3860) : 0
(95152,3440):(95372,3860) : 1
(95152,3440):(95372,3860) : 2
(95152,3440):(95372,3860) : 3
D[13]
use : s
dir : i
shape : 
(97316,3440):(97536,3860) : 0
(97316,3440):(97536,3860) : 1
(97316,3440):(97536,3860) : 2
(97316,3440):(97536,3860) : 3
D[14]
use : s
dir : i
shape : 
(107288,3440):(107508,3860) : 0
(107288,3440):(107508,3860) : 1
(107288,3440):(107508,3860) : 2
(107288,3440):(107508,3860) : 3
D[15]
use : s
dir : i
shape : 
(109452,3440):(109672,3860) : 0
(109452,3440):(109672,3860) : 1
(109452,3440):(109672,3860) : 2
(109452,3440):(109672,3860) : 3
D[1]
use : s
dir : i
shape : 
(11256,3440):(11476,3860) : 0
(11256,3440):(11476,3860) : 1
(11256,3440):(11476,3860) : 2
(11256,3440):(11476,3860) : 3
D[2]
use : s
dir : i
shape : 
(21228,3440):(21448,3860) : 0
(21228,3440):(21448,3860) : 1
(21228,3440):(21448,3860) : 2
(21228,3440):(21448,3860) : 3
D[3]
use : s
dir : i
shape : 
(23392,3440):(23612,3860) : 0
(23392,3440):(23612,3860) : 1
(23392,3440):(23612,3860) : 2
(23392,3440):(23612,3860) : 3
D[4]
use : s
dir : i
shape : 
(33364,3440):(33584,3860) : 0
(33364,3440):(33584,3860) : 1
(33364,3440):(33584,3860) : 2
(33364,3440):(33584,3860) : 3
D[5]
use : s
dir : i
shape : 
(35528,3440):(35748,3860) : 0
(35528,3440):(35748,3860) : 1
(35528,3440):(35748,3860) : 2
(35528,3440):(35748,3860) : 3
D[6]
use : s
dir : i
shape : 
(45500,3440):(45720,3860) : 0
(45500,3440):(45720,3860) : 1
(45500,3440):(45720,3860) : 2
(45500,3440):(45720,3860) : 3
D[7]
use : s
dir : i
shape : 
(47664,3440):(47884,3860) : 0
(47664,3440):(47884,3860) : 1
(47664,3440):(47884,3860) : 2
(47664,3440):(47884,3860) : 3
D[8]
use : s
dir : i
shape : 
(70880,3440):(71100,3860) : 0
(70880,3440):(71100,3860) : 1
(70880,3440):(71100,3860) : 2
(70880,3440):(71100,3860) : 3
D[9]
use : s
dir : i
shape : 
(73044,3440):(73264,3860) : 0
(73044,3440):(73264,3860) : 1
(73044,3440):(73264,3860) : 2
(73044,3440):(73264,3860) : 3
OEN
use : s
dir : i
shape : 
(65160,3440):(65380,3860) : 0
(65160,3440):(65380,3860) : 1
(65160,3440):(65380,3860) : 2
(65160,3440):(65380,3860) : 3
Q[0]
use : s
dir :  
shape : 
(7996,3440):(8216,3860) : 0
(7996,3440):(8216,3860) : 1
(7996,3440):(8216,3860) : 2
(7996,3440):(8216,3860) : 3
Q[10]
use : s
dir :  
shape : 
(81960,3440):(82180,3860) : 0
(81960,3440):(82180,3860) : 1
(81960,3440):(82180,3860) : 2
(81960,3440):(82180,3860) : 3
Q[11]
use : s
dir :  
shape : 
(86236,3440):(86456,3860) : 0
(86236,3440):(86456,3860) : 1
(86236,3440):(86456,3860) : 2
(86236,3440):(86456,3860) : 3
Q[12]
use : s
dir :  
shape : 
(94096,3440):(94316,3860) : 0
(94096,3440):(94316,3860) : 1
(94096,3440):(94316,3860) : 2
(94096,3440):(94316,3860) : 3
Q[13]
use : s
dir :  
shape : 
(98372,3440):(98592,3860) : 0
(98372,3440):(98592,3860) : 1
(98372,3440):(98592,3860) : 2
(98372,3440):(98592,3860) : 3
Q[14]
use : s
dir :  
shape : 
(106232,3440):(106452,3860) : 0
(106232,3440):(106452,3860) : 1
(106232,3440):(106452,3860) : 2
(106232,3440):(106452,3860) : 3
Q[15]
use : s
dir :  
shape : 
(110528,3440):(110748,3860) : 0
(110528,3440):(110748,3860) : 1
(110528,3440):(110748,3860) : 2
(110528,3440):(110748,3860) : 3
Q[1]
use : s
dir :  
shape : 
(12312,3440):(12532,3860) : 0
(12312,3440):(12532,3860) : 1
(12312,3440):(12532,3860) : 2
(12312,3440):(12532,3860) : 3
Q[2]
use : s
dir :  
shape : 
(20172,3440):(20392,3860) : 0
(20172,3440):(20392,3860) : 1
(20172,3440):(20392,3860) : 2
(20172,3440):(20392,3860) : 3
Q[3]
use : s
dir :  
shape : 
(24448,3440):(24668,3860) : 0
(24448,3440):(24668,3860) : 1
(24448,3440):(24668,3860) : 2
(24448,3440):(24668,3860) : 3
Q[4]
use : s
dir :  
shape : 
(32308,3440):(32528,3860) : 0
(32308,3440):(32528,3860) : 1
(32308,3440):(32528,3860) : 2
(32308,3440):(32528,3860) : 3
Q[5]
use : s
dir :  
shape : 
(36584,3440):(36804,3860) : 0
(36584,3440):(36804,3860) : 1
(36584,3440):(36804,3860) : 2
(36584,3440):(36804,3860) : 3
Q[6]
use : s
dir :  
shape : 
(44444,3440):(44664,3860) : 0
(44444,3440):(44664,3860) : 1
(44444,3440):(44664,3860) : 2
(44444,3440):(44664,3860) : 3
Q[7]
use : s
dir :  
shape : 
(48720,3440):(48940,3860) : 0
(48720,3440):(48940,3860) : 1
(48720,3440):(48940,3860) : 2
(48720,3440):(48940,3860) : 3
Q[8]
use : s
dir :  
shape : 
(69824,3440):(70044,3860) : 0
(69824,3440):(70044,3860) : 1
(69824,3440):(70044,3860) : 2
(69824,3440):(70044,3860) : 3
Q[9]
use : s
dir :  
shape : 
(74100,3440):(74320,3860) : 0
(74100,3440):(74320,3860) : 1
(74100,3440):(74320,3860) : 2
(74100,3440):(74320,3860) : 3
WEN
use : s
dir : i
shape : 
(63432,3440):(63652,3860) : 0
(63432,3440):(63652,3860) : 1
(63432,3440):(63652,3860) : 2
(63432,3440):(63652,3860) : 3
VDD
use : p
dir : b
shape : 
(0,32400):(118764,33800) : 4
(0,0):(118764,1400) : 4
(117364,0):(118764,33798) : 3
(0,0):(1400,33798) : 3
VSS
use : g
dir : b
shape : 
(1720,30680):(117044,32080) : 4
(1720,1720):(117044,3120) : 4
(115644,1720):(117044,32080) : 3
(1720,1720):(3120,32080) : 3
PCORNERDG
--pins(0)
PDIDGZ
--pins(2)
PAD
use :  
dir : i
shape : 
(3754,0):(4448,272) : 0
(3754,0):(4448,272) : 1
C
use :  
dir : o
shape : 
(6434,46800):(6834,47000) : 0
(6434,46800):(6834,47000) : 1
(6434,46800):(6834,47000) : 2
(6434,46800):(6834,47000) : 3
(6434,46800):(6834,47000) : 4
PDO04CDG
--pins(2)
PAD
use :  
dir : o
shape : 
(3754,0):(4448,272) : 0
(3754,0):(4448,272) : 1
I
use :  
dir : i
shape : 
(6434,46800):(6834,47000) : 0
(6434,46800):(6834,47000) : 1
(6434,46800):(6834,47000) : 2
(6434,46800):(6834,47000) : 3
(6434,46800):(6834,47000) : 4
PVDD1DGZ
--pins(1)
VDD
use : p
dir : o
shape : 
(1200,45400):(6800,47000) : 2
(1200,45400):(6800,47000) : 3
(1200,45400):(6800,47000) : 4
PVSS1DGZ
--pins(1)
VSS
use : g
dir : o
shape : 
(1200,45400):(6800,47000) : 2
(1200,45400):(6800,47000) : 3
(1200,45400):(6800,47000) : 4
Metal1 (V) p200,200 w100 s120 a46000 prefer: srt100 stp200 num1953 wrong: srt200 stp200 num1949
Metal2 (H) p200,200 w100 s160 a56000 prefer: srt200 stp200 num1949 wrong: srt100 stp200 num1953
Metal3 (V) p200,200 w100 s160 a68000 prefer: srt100 stp200 num1953 wrong: srt200 stp200 num1949
Metal4 (H) p200,200 w100 s160 a68000 prefer: srt200 stp200 num1949 wrong: srt100 stp200 num1953
Metal5 (V) p200,200 w100 s160 a68000 prefer: srt100 stp200 num1953 wrong: srt200 stp200 num1949
Metal6 (H) p300,300 w140 s200 a100000 prefer: srt200 stp300 num1300 wrong: srt400 stp300 num1301
Metal7 (V) p300,300 w140 s200 a100000 prefer: srt400 stp300 num1301 wrong: srt200 stp300 num1300
Metal8 (H) p400,400 w200 s240 a208000 prefer: srt200 stp400 num975 wrong: srt500 stp400 num976
Metal9 (V) p400,400 w200 s240 a208000 prefer: srt500 stp400 num976 wrong: srt200 stp400 num975
